LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY LGC_Netlist IS
    PORT (
        clk : IN STD_LOGIC;
        rst : IN STD_LOGIC;
        readyMEM : IN STD_LOGIC;
        dataBusIn : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
        p1TRF : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
        p2TRF : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		PbarS : IN STD_LOGIC;				-- added for scan insertion
		Si_3 : IN STD_LOGIC;                -- added for scan insertion
		Si_4 : IN STD_LOGIC;                -- added for scan insertion
		Si_5 : IN STD_LOGIC;                -- added for scan insertion
		Si_6 : IN STD_LOGIC;                -- added for scan insertion
		So_1 : OUT STD_LOGIC;               -- added for scan insertion
		So_2 : OUT STD_LOGIC;               -- added for scan insertion
		So_3 : OUT STD_LOGIC;               -- added for scan insertion
		So_4 : OUT STD_LOGIC;               -- added for scan insertion
		readMM : OUT STD_LOGIC;
        writeMM : OUT STD_LOGIC;
        dataBusOut : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
        addrBus : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
        outMuxrs1 : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
        outMuxrs2 : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
        outMuxrd : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
        inDataTRF : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
        writeTRF : OUT STD_LOGIC;
        readInst : OUT STD_LOGIC);
END ENTITY LGC_Netlist;

ARCHITECTURE arch OF LGC_Netlist IS
    SIGNAL PbarS_sig : STD_LOGIC;		                    -- added for scan insertion
	SIGNAL Si_3_sig : STD_LOGIC;                            -- added for scan insertion
	SIGNAL Si_4_sig : STD_LOGIC;                            -- added for scan insertion
	SIGNAL Si_5_sig : STD_LOGIC;                            -- added for scan insertion
	SIGNAL Si_6_sig : STD_LOGIC;                            -- added for scan insertion
	SIGNAL So_1_sig : STD_LOGIC;                            -- added for scan insertion
	SIGNAL So_2_sig : STD_LOGIC;                            -- added for scan insertion
	SIGNAL So_3_sig : STD_LOGIC;                            -- added for scan insertion
	SIGNAL So_4_sig : STD_LOGIC;                            -- added for scan insertion
    SIGNAL fakeDFF_sig : STD_LOGIC_VECTOR (9 DOWNTO 0);    -- added for scan insertion
	
	SIGNAL S0 : STD_LOGIC;
    SIGNAL S1 : STD_LOGIC;
    SIGNAL S2 : STD_LOGIC;
    SIGNAL S3 : STD_LOGIC;
    SIGNAL S4 : STD_LOGIC;
    SIGNAL S5 : STD_LOGIC;
    SIGNAL S6 : STD_LOGIC;
    SIGNAL S7 : STD_LOGIC;
    SIGNAL S8 : STD_LOGIC;
    SIGNAL S9 : STD_LOGIC;
    SIGNAL S10 : STD_LOGIC;
    SIGNAL S11 : STD_LOGIC;
    SIGNAL S12 : STD_LOGIC;
    SIGNAL S13 : STD_LOGIC;
    SIGNAL S14 : STD_LOGIC;
    SIGNAL S15 : STD_LOGIC;
    SIGNAL S16 : STD_LOGIC;
    SIGNAL S17 : STD_LOGIC;
    SIGNAL S18 : STD_LOGIC;
    SIGNAL S19 : STD_LOGIC;
    SIGNAL S20 : STD_LOGIC;
    SIGNAL S21 : STD_LOGIC;
    SIGNAL S22 : STD_LOGIC;
    SIGNAL S23 : STD_LOGIC;
    SIGNAL S24 : STD_LOGIC;
    SIGNAL S25 : STD_LOGIC;
    SIGNAL S26 : STD_LOGIC;
    SIGNAL S27 : STD_LOGIC;
    SIGNAL S28 : STD_LOGIC;
    SIGNAL S29 : STD_LOGIC;
    SIGNAL S30 : STD_LOGIC;
    SIGNAL S31 : STD_LOGIC;
    SIGNAL S32 : STD_LOGIC;
    SIGNAL S33 : STD_LOGIC;
    SIGNAL S34 : STD_LOGIC;
    SIGNAL S35 : STD_LOGIC;
    SIGNAL S36 : STD_LOGIC;
    SIGNAL S37 : STD_LOGIC;
    SIGNAL S38 : STD_LOGIC;
    SIGNAL S39 : STD_LOGIC;
    SIGNAL S40 : STD_LOGIC;
    SIGNAL S41 : STD_LOGIC;
    SIGNAL S42 : STD_LOGIC;
    SIGNAL S43 : STD_LOGIC;
    SIGNAL S44 : STD_LOGIC;
    SIGNAL S45 : STD_LOGIC;
    SIGNAL S46 : STD_LOGIC;
    SIGNAL S47 : STD_LOGIC;
    SIGNAL S48 : STD_LOGIC;
    SIGNAL S49 : STD_LOGIC;
    SIGNAL S50 : STD_LOGIC;
    SIGNAL S51 : STD_LOGIC;
    SIGNAL S52 : STD_LOGIC;
    SIGNAL S53 : STD_LOGIC;
    SIGNAL S54 : STD_LOGIC;
    SIGNAL S55 : STD_LOGIC;
    SIGNAL S56 : STD_LOGIC;
    SIGNAL S57 : STD_LOGIC;
    SIGNAL S58 : STD_LOGIC;
    SIGNAL S59 : STD_LOGIC;
    SIGNAL S60 : STD_LOGIC;
    SIGNAL S61 : STD_LOGIC;
    SIGNAL S62 : STD_LOGIC;
    SIGNAL S63 : STD_LOGIC;
    SIGNAL S64 : STD_LOGIC;
    SIGNAL S65 : STD_LOGIC;
    SIGNAL S66 : STD_LOGIC;
    SIGNAL S67 : STD_LOGIC;
    SIGNAL S68 : STD_LOGIC;
    SIGNAL S69 : STD_LOGIC;
    SIGNAL S70 : STD_LOGIC;
    SIGNAL S71 : STD_LOGIC;
    SIGNAL S72 : STD_LOGIC;
    SIGNAL S73 : STD_LOGIC;
    SIGNAL S74 : STD_LOGIC;
    SIGNAL S75 : STD_LOGIC;
    SIGNAL S76 : STD_LOGIC;
    SIGNAL S77 : STD_LOGIC;
    SIGNAL S78 : STD_LOGIC;
    SIGNAL S79 : STD_LOGIC;
    SIGNAL S80 : STD_LOGIC;
    SIGNAL S81 : STD_LOGIC;
    SIGNAL S82 : STD_LOGIC;
    SIGNAL S83 : STD_LOGIC;
    SIGNAL S84 : STD_LOGIC;
    SIGNAL S85 : STD_LOGIC;
    SIGNAL S86 : STD_LOGIC;
    SIGNAL S87 : STD_LOGIC;
    SIGNAL S88 : STD_LOGIC;
    SIGNAL S89 : STD_LOGIC;
    SIGNAL S90 : STD_LOGIC;
    SIGNAL S91 : STD_LOGIC;
    SIGNAL S92 : STD_LOGIC;
    SIGNAL S93 : STD_LOGIC;
    SIGNAL S94 : STD_LOGIC;
    SIGNAL S95 : STD_LOGIC;
    SIGNAL S96 : STD_LOGIC;
    SIGNAL S97 : STD_LOGIC;
    SIGNAL S98 : STD_LOGIC;
    SIGNAL S99 : STD_LOGIC;
    SIGNAL S100 : STD_LOGIC;
    SIGNAL S101 : STD_LOGIC;
    SIGNAL S102 : STD_LOGIC;
    SIGNAL S103 : STD_LOGIC;
    SIGNAL S104 : STD_LOGIC;
    SIGNAL S105 : STD_LOGIC;
    SIGNAL S106 : STD_LOGIC;
    SIGNAL S107 : STD_LOGIC;
    SIGNAL S108 : STD_LOGIC;
    SIGNAL S109 : STD_LOGIC;
    SIGNAL S110 : STD_LOGIC;
    SIGNAL S111 : STD_LOGIC;
    SIGNAL S112 : STD_LOGIC;
    SIGNAL S113 : STD_LOGIC;
    SIGNAL S114 : STD_LOGIC;
    SIGNAL S115 : STD_LOGIC;
    SIGNAL S116 : STD_LOGIC;
    SIGNAL S117 : STD_LOGIC;
    SIGNAL S118 : STD_LOGIC;
    SIGNAL S119 : STD_LOGIC;
    SIGNAL S120 : STD_LOGIC;
    SIGNAL S121 : STD_LOGIC;
    SIGNAL S122 : STD_LOGIC;
    SIGNAL S123 : STD_LOGIC;
    SIGNAL S124 : STD_LOGIC;
    SIGNAL S125 : STD_LOGIC;
    SIGNAL S126 : STD_LOGIC;
    SIGNAL S127 : STD_LOGIC;
    SIGNAL S128 : STD_LOGIC;
    SIGNAL S129 : STD_LOGIC;
    SIGNAL S130 : STD_LOGIC;
    SIGNAL S131 : STD_LOGIC;
    SIGNAL S132 : STD_LOGIC;
    SIGNAL S133 : STD_LOGIC;
    SIGNAL S134 : STD_LOGIC;
    SIGNAL S135 : STD_LOGIC;
    SIGNAL S136 : STD_LOGIC;
    SIGNAL S137 : STD_LOGIC;
    SIGNAL S138 : STD_LOGIC;
    SIGNAL S139 : STD_LOGIC;
    SIGNAL S140 : STD_LOGIC;
    SIGNAL S141 : STD_LOGIC;
    SIGNAL S142 : STD_LOGIC;
    SIGNAL S143 : STD_LOGIC;
    SIGNAL S144 : STD_LOGIC;
    SIGNAL S145 : STD_LOGIC;
    SIGNAL S146 : STD_LOGIC;
    SIGNAL S147 : STD_LOGIC;
    SIGNAL S148 : STD_LOGIC;
    SIGNAL S149 : STD_LOGIC;
    SIGNAL S150 : STD_LOGIC;
    SIGNAL S151 : STD_LOGIC;
    SIGNAL S152 : STD_LOGIC;
    SIGNAL S153 : STD_LOGIC;
    SIGNAL S154 : STD_LOGIC;
    SIGNAL S155 : STD_LOGIC;
    SIGNAL S156 : STD_LOGIC;
    SIGNAL S157 : STD_LOGIC;
    SIGNAL S158 : STD_LOGIC;
    SIGNAL S159 : STD_LOGIC;
    SIGNAL S160 : STD_LOGIC;
    SIGNAL S161 : STD_LOGIC;
    SIGNAL S162 : STD_LOGIC;
    SIGNAL S163 : STD_LOGIC;
    SIGNAL S164 : STD_LOGIC;
    SIGNAL S165 : STD_LOGIC;
    SIGNAL S166 : STD_LOGIC;
    SIGNAL S167 : STD_LOGIC;
    SIGNAL S168 : STD_LOGIC;
    SIGNAL S169 : STD_LOGIC;
    SIGNAL S170 : STD_LOGIC;
    SIGNAL S171 : STD_LOGIC;
    SIGNAL S172 : STD_LOGIC;
    SIGNAL S173 : STD_LOGIC;
    SIGNAL S174 : STD_LOGIC;
    SIGNAL S175 : STD_LOGIC;
    SIGNAL S176 : STD_LOGIC;
    SIGNAL S177 : STD_LOGIC;
    SIGNAL S178 : STD_LOGIC;
    SIGNAL S179 : STD_LOGIC;
    SIGNAL S180 : STD_LOGIC;
    SIGNAL S181 : STD_LOGIC;
    SIGNAL S182 : STD_LOGIC;
    SIGNAL S183 : STD_LOGIC;
    SIGNAL S184 : STD_LOGIC;
    SIGNAL S185 : STD_LOGIC;
    SIGNAL S186 : STD_LOGIC;
    SIGNAL S187 : STD_LOGIC;
    SIGNAL S188 : STD_LOGIC;
    SIGNAL S189 : STD_LOGIC;
    SIGNAL S190 : STD_LOGIC;
    SIGNAL S191 : STD_LOGIC;
    SIGNAL S192 : STD_LOGIC;
    SIGNAL S193 : STD_LOGIC;
    SIGNAL S194 : STD_LOGIC;
    SIGNAL S195 : STD_LOGIC;
    SIGNAL S196 : STD_LOGIC;
    SIGNAL S197 : STD_LOGIC;
    SIGNAL S198 : STD_LOGIC;
    SIGNAL S199 : STD_LOGIC;
    SIGNAL S200 : STD_LOGIC;
    SIGNAL S201 : STD_LOGIC;
    SIGNAL S202 : STD_LOGIC;
    SIGNAL S203 : STD_LOGIC;
    SIGNAL S204 : STD_LOGIC;
    SIGNAL S205 : STD_LOGIC;
    SIGNAL S206 : STD_LOGIC;
    SIGNAL S207 : STD_LOGIC;
    SIGNAL S208 : STD_LOGIC;
    SIGNAL S209 : STD_LOGIC;
    SIGNAL S210 : STD_LOGIC;
    SIGNAL S211 : STD_LOGIC;
    SIGNAL S212 : STD_LOGIC;
    SIGNAL S213 : STD_LOGIC;
    SIGNAL S214 : STD_LOGIC;
    SIGNAL S215 : STD_LOGIC;
    SIGNAL S216 : STD_LOGIC;
    SIGNAL S217 : STD_LOGIC;
    SIGNAL S218 : STD_LOGIC;
    SIGNAL S219 : STD_LOGIC;
    SIGNAL S220 : STD_LOGIC;
    SIGNAL S221 : STD_LOGIC;
    SIGNAL S222 : STD_LOGIC;
    SIGNAL S223 : STD_LOGIC;
    SIGNAL S224 : STD_LOGIC;
    SIGNAL S225 : STD_LOGIC;
    SIGNAL S226 : STD_LOGIC;
    SIGNAL S227 : STD_LOGIC;
    SIGNAL S228 : STD_LOGIC;
    SIGNAL S229 : STD_LOGIC;
    SIGNAL S230 : STD_LOGIC;
    SIGNAL S231 : STD_LOGIC;
    SIGNAL S232 : STD_LOGIC;
    SIGNAL S233 : STD_LOGIC;
    SIGNAL S234 : STD_LOGIC;
    SIGNAL S235 : STD_LOGIC;
    SIGNAL S236 : STD_LOGIC;
    SIGNAL S237 : STD_LOGIC;
    SIGNAL S238 : STD_LOGIC;
    SIGNAL S239 : STD_LOGIC;
    SIGNAL S240 : STD_LOGIC;
    SIGNAL S241 : STD_LOGIC;
    SIGNAL S242 : STD_LOGIC;
    SIGNAL S243 : STD_LOGIC;
    SIGNAL S244 : STD_LOGIC;
    SIGNAL S245 : STD_LOGIC;
    SIGNAL S246 : STD_LOGIC;
    SIGNAL S247 : STD_LOGIC;
    SIGNAL S248 : STD_LOGIC;
    SIGNAL S249 : STD_LOGIC;
    SIGNAL S250 : STD_LOGIC;
    SIGNAL S251 : STD_LOGIC;
    SIGNAL S252 : STD_LOGIC;
    SIGNAL S253 : STD_LOGIC;
    SIGNAL S254 : STD_LOGIC;
    SIGNAL S255 : STD_LOGIC;
    SIGNAL S256 : STD_LOGIC;
    SIGNAL S257 : STD_LOGIC;
    SIGNAL S258 : STD_LOGIC;
    SIGNAL S259 : STD_LOGIC;
    SIGNAL S260 : STD_LOGIC;
    SIGNAL S261 : STD_LOGIC;
    SIGNAL S262 : STD_LOGIC;
    SIGNAL S263 : STD_LOGIC;
    SIGNAL S264 : STD_LOGIC;
    SIGNAL S265 : STD_LOGIC;
    SIGNAL S266 : STD_LOGIC;
    SIGNAL S267 : STD_LOGIC;
    SIGNAL S268 : STD_LOGIC;
    SIGNAL S269 : STD_LOGIC;
    SIGNAL S270 : STD_LOGIC;
    SIGNAL S271 : STD_LOGIC;
    SIGNAL S272 : STD_LOGIC;
    SIGNAL S273 : STD_LOGIC;
    SIGNAL S274 : STD_LOGIC;
    SIGNAL S275 : STD_LOGIC;
    SIGNAL S276 : STD_LOGIC;
    SIGNAL S277 : STD_LOGIC;
    SIGNAL S278 : STD_LOGIC;
    SIGNAL S279 : STD_LOGIC;
    SIGNAL S280 : STD_LOGIC;
    SIGNAL S281 : STD_LOGIC;
    SIGNAL S282 : STD_LOGIC;
    SIGNAL S283 : STD_LOGIC;
    SIGNAL S284 : STD_LOGIC;
    SIGNAL S285 : STD_LOGIC;
    SIGNAL S286 : STD_LOGIC;
    SIGNAL S287 : STD_LOGIC;
    SIGNAL S288 : STD_LOGIC;
    SIGNAL S289 : STD_LOGIC;
    SIGNAL S290 : STD_LOGIC;
    SIGNAL S291 : STD_LOGIC;
    SIGNAL S292 : STD_LOGIC;
    SIGNAL S293 : STD_LOGIC;
    SIGNAL S294 : STD_LOGIC;
    SIGNAL S295 : STD_LOGIC;
    SIGNAL S296 : STD_LOGIC;
    SIGNAL S297 : STD_LOGIC;
    SIGNAL S298 : STD_LOGIC;
    SIGNAL S299 : STD_LOGIC;
    SIGNAL S300 : STD_LOGIC;
    SIGNAL S301 : STD_LOGIC;
    SIGNAL S302 : STD_LOGIC;
    SIGNAL S303 : STD_LOGIC;
    SIGNAL S304 : STD_LOGIC;
    SIGNAL S305 : STD_LOGIC;
    SIGNAL S306 : STD_LOGIC;
    SIGNAL S307 : STD_LOGIC;
    SIGNAL S308 : STD_LOGIC;
    SIGNAL S309 : STD_LOGIC;
    SIGNAL S310 : STD_LOGIC;
    SIGNAL S311 : STD_LOGIC;
    SIGNAL S312 : STD_LOGIC;
    SIGNAL S313 : STD_LOGIC;
    SIGNAL S314 : STD_LOGIC;
    SIGNAL S315 : STD_LOGIC;
    SIGNAL S316 : STD_LOGIC;
    SIGNAL S317 : STD_LOGIC;
    SIGNAL S318 : STD_LOGIC;
    SIGNAL S319 : STD_LOGIC;
    SIGNAL S320 : STD_LOGIC;
    SIGNAL S321 : STD_LOGIC;
    SIGNAL S322 : STD_LOGIC;
    SIGNAL S323 : STD_LOGIC;
    SIGNAL S324 : STD_LOGIC;
    SIGNAL S325 : STD_LOGIC;
    SIGNAL S326 : STD_LOGIC;
    SIGNAL S327 : STD_LOGIC;
    SIGNAL S328 : STD_LOGIC;
    SIGNAL S329 : STD_LOGIC;
    SIGNAL S330 : STD_LOGIC;
    SIGNAL S331 : STD_LOGIC;
    SIGNAL S332 : STD_LOGIC;
    SIGNAL S333 : STD_LOGIC;
    SIGNAL S334 : STD_LOGIC;
    SIGNAL S335 : STD_LOGIC;
    SIGNAL S336 : STD_LOGIC;
    SIGNAL S337 : STD_LOGIC;
    SIGNAL S338 : STD_LOGIC;
    SIGNAL S339 : STD_LOGIC;
    SIGNAL S340 : STD_LOGIC;
    SIGNAL S341 : STD_LOGIC;
    SIGNAL S342 : STD_LOGIC;
    SIGNAL S343 : STD_LOGIC;
    SIGNAL S344 : STD_LOGIC;
    SIGNAL S345 : STD_LOGIC;
    SIGNAL S346 : STD_LOGIC;
    SIGNAL S347 : STD_LOGIC;
    SIGNAL S348 : STD_LOGIC;
    SIGNAL S349 : STD_LOGIC;
    SIGNAL S350 : STD_LOGIC;
    SIGNAL S351 : STD_LOGIC;
    SIGNAL S352 : STD_LOGIC;
    SIGNAL S353 : STD_LOGIC;
    SIGNAL S354 : STD_LOGIC;
    SIGNAL S355 : STD_LOGIC;
    SIGNAL S356 : STD_LOGIC;
    SIGNAL S357 : STD_LOGIC;
    SIGNAL S358 : STD_LOGIC;
    SIGNAL S359 : STD_LOGIC;
    SIGNAL S360 : STD_LOGIC;
    SIGNAL S361 : STD_LOGIC;
    SIGNAL S362 : STD_LOGIC;
    SIGNAL S363 : STD_LOGIC;
    SIGNAL S364 : STD_LOGIC;
    SIGNAL S365 : STD_LOGIC;
    SIGNAL S366 : STD_LOGIC;
    SIGNAL S367 : STD_LOGIC;
    SIGNAL S368 : STD_LOGIC;
    SIGNAL S369 : STD_LOGIC;
    SIGNAL S370 : STD_LOGIC;
    SIGNAL S371 : STD_LOGIC;
    SIGNAL S372 : STD_LOGIC;
    SIGNAL S373 : STD_LOGIC;
    SIGNAL S374 : STD_LOGIC;
    SIGNAL S375 : STD_LOGIC;
    SIGNAL S376 : STD_LOGIC;
    SIGNAL S377 : STD_LOGIC;
    SIGNAL S378 : STD_LOGIC;
    SIGNAL S379 : STD_LOGIC;
    SIGNAL S380 : STD_LOGIC;
    SIGNAL S381 : STD_LOGIC;
    SIGNAL S382 : STD_LOGIC;
    SIGNAL S383 : STD_LOGIC;
    SIGNAL S384 : STD_LOGIC;
    SIGNAL S385 : STD_LOGIC;
    SIGNAL S386 : STD_LOGIC;
    SIGNAL S387 : STD_LOGIC;
    SIGNAL S388 : STD_LOGIC;
    SIGNAL S389 : STD_LOGIC;
    SIGNAL S390 : STD_LOGIC;
    SIGNAL S391 : STD_LOGIC;
    SIGNAL S392 : STD_LOGIC;
    SIGNAL S393 : STD_LOGIC;
    SIGNAL S394 : STD_LOGIC;
    SIGNAL S395 : STD_LOGIC;
    SIGNAL S396 : STD_LOGIC;
    SIGNAL S397 : STD_LOGIC;
    SIGNAL S398 : STD_LOGIC;
    SIGNAL S399 : STD_LOGIC;
    SIGNAL S400 : STD_LOGIC;
    SIGNAL S401 : STD_LOGIC;
    SIGNAL S402 : STD_LOGIC;
    SIGNAL S403 : STD_LOGIC;
    SIGNAL S404 : STD_LOGIC;
    SIGNAL S405 : STD_LOGIC;
    SIGNAL S406 : STD_LOGIC;
    SIGNAL S407 : STD_LOGIC;
    SIGNAL S408 : STD_LOGIC;
    SIGNAL S409 : STD_LOGIC;
    SIGNAL S410 : STD_LOGIC;
    SIGNAL S411 : STD_LOGIC;
    SIGNAL S412 : STD_LOGIC;
    SIGNAL S413 : STD_LOGIC;
    SIGNAL S414 : STD_LOGIC;
    SIGNAL S415 : STD_LOGIC;
    SIGNAL S416 : STD_LOGIC;
    SIGNAL S417 : STD_LOGIC;
    SIGNAL S418 : STD_LOGIC;
    SIGNAL S419 : STD_LOGIC;
    SIGNAL S420 : STD_LOGIC;
    SIGNAL S421 : STD_LOGIC;
    SIGNAL S422 : STD_LOGIC;
    SIGNAL S423 : STD_LOGIC;
    SIGNAL S424 : STD_LOGIC;
    SIGNAL S425 : STD_LOGIC;
    SIGNAL S426 : STD_LOGIC;
    SIGNAL S427 : STD_LOGIC;
    SIGNAL S428 : STD_LOGIC;
    SIGNAL S429 : STD_LOGIC;
    SIGNAL S430 : STD_LOGIC;
    SIGNAL S431 : STD_LOGIC;
    SIGNAL S432 : STD_LOGIC;
    SIGNAL S433 : STD_LOGIC;
    SIGNAL S434 : STD_LOGIC;
    SIGNAL S435 : STD_LOGIC;
    SIGNAL S436 : STD_LOGIC;
    SIGNAL S437 : STD_LOGIC;
    SIGNAL S438 : STD_LOGIC;
    SIGNAL S439 : STD_LOGIC;
    SIGNAL S440 : STD_LOGIC;
    SIGNAL S441 : STD_LOGIC;
    SIGNAL S442 : STD_LOGIC;
    SIGNAL S443 : STD_LOGIC;
    SIGNAL S444 : STD_LOGIC;
    SIGNAL S445 : STD_LOGIC;
    SIGNAL S446 : STD_LOGIC;
    SIGNAL S447 : STD_LOGIC;
    SIGNAL S448 : STD_LOGIC;
    SIGNAL S449 : STD_LOGIC;
    SIGNAL S450 : STD_LOGIC;
    SIGNAL S451 : STD_LOGIC;
    SIGNAL S452 : STD_LOGIC;
    SIGNAL S453 : STD_LOGIC;
    SIGNAL S454 : STD_LOGIC;
    SIGNAL S455 : STD_LOGIC;
    SIGNAL S456 : STD_LOGIC;
    SIGNAL S457 : STD_LOGIC;
    SIGNAL S458 : STD_LOGIC;
    SIGNAL S459 : STD_LOGIC;
    SIGNAL S460 : STD_LOGIC;
    SIGNAL S461 : STD_LOGIC;
    SIGNAL S462 : STD_LOGIC;
    SIGNAL S463 : STD_LOGIC;
    SIGNAL S464 : STD_LOGIC;
    SIGNAL S465 : STD_LOGIC;
    SIGNAL S466 : STD_LOGIC;
    SIGNAL S467 : STD_LOGIC;
    SIGNAL S468 : STD_LOGIC;
    SIGNAL S469 : STD_LOGIC;
    SIGNAL S470 : STD_LOGIC;
    SIGNAL S471 : STD_LOGIC;
    SIGNAL S472 : STD_LOGIC;
    SIGNAL S473 : STD_LOGIC;
    SIGNAL S474 : STD_LOGIC;
    SIGNAL S475 : STD_LOGIC;
    SIGNAL S476 : STD_LOGIC;
    SIGNAL S477 : STD_LOGIC;
    SIGNAL S478 : STD_LOGIC;
    SIGNAL S479 : STD_LOGIC;
    SIGNAL S480 : STD_LOGIC;
    SIGNAL S481 : STD_LOGIC;
    SIGNAL S482 : STD_LOGIC;
    SIGNAL S483 : STD_LOGIC;
    SIGNAL S484 : STD_LOGIC;
    SIGNAL S485 : STD_LOGIC;
    SIGNAL S486 : STD_LOGIC;
    SIGNAL S487 : STD_LOGIC;
    SIGNAL S488 : STD_LOGIC;
    SIGNAL S489 : STD_LOGIC;
    SIGNAL S490 : STD_LOGIC;
    SIGNAL S491 : STD_LOGIC;
    SIGNAL S492 : STD_LOGIC;
    SIGNAL S493 : STD_LOGIC;
    SIGNAL S494 : STD_LOGIC;
    SIGNAL S495 : STD_LOGIC;
    SIGNAL S496 : STD_LOGIC;
    SIGNAL S497 : STD_LOGIC;
    SIGNAL S498 : STD_LOGIC;
    SIGNAL S499 : STD_LOGIC;
    SIGNAL S500 : STD_LOGIC;
    SIGNAL S501 : STD_LOGIC;
    SIGNAL S502 : STD_LOGIC;
    SIGNAL S503 : STD_LOGIC;
    SIGNAL S504 : STD_LOGIC;
    SIGNAL S505 : STD_LOGIC;
    SIGNAL S506 : STD_LOGIC;
    SIGNAL S507 : STD_LOGIC;
    SIGNAL S508 : STD_LOGIC;
    SIGNAL S509 : STD_LOGIC;
    SIGNAL S510 : STD_LOGIC;
    SIGNAL S511 : STD_LOGIC;
    SIGNAL S512 : STD_LOGIC;
    SIGNAL S513 : STD_LOGIC;
    SIGNAL S514 : STD_LOGIC;
    SIGNAL S515 : STD_LOGIC;
    SIGNAL S516 : STD_LOGIC;
    SIGNAL S517 : STD_LOGIC;
    SIGNAL S518 : STD_LOGIC;
    SIGNAL S519 : STD_LOGIC;
    SIGNAL S520 : STD_LOGIC;
    SIGNAL S521 : STD_LOGIC;
    SIGNAL S522 : STD_LOGIC;
    SIGNAL S523 : STD_LOGIC;
    SIGNAL S524 : STD_LOGIC;
    SIGNAL S525 : STD_LOGIC;
    SIGNAL S526 : STD_LOGIC;
    SIGNAL S527 : STD_LOGIC;
    SIGNAL S528 : STD_LOGIC;
    SIGNAL S529 : STD_LOGIC;
    SIGNAL S530 : STD_LOGIC;
    SIGNAL S531 : STD_LOGIC;
    SIGNAL S532 : STD_LOGIC;
    SIGNAL S533 : STD_LOGIC;
    SIGNAL S534 : STD_LOGIC;
    SIGNAL S535 : STD_LOGIC;
    SIGNAL S536 : STD_LOGIC;
    SIGNAL S537 : STD_LOGIC;
    SIGNAL S538 : STD_LOGIC;
    SIGNAL S539 : STD_LOGIC;
    SIGNAL S540 : STD_LOGIC;
    SIGNAL S541 : STD_LOGIC;
    SIGNAL S542 : STD_LOGIC;
    SIGNAL S543 : STD_LOGIC;
    SIGNAL S544 : STD_LOGIC;
    SIGNAL S545 : STD_LOGIC;
    SIGNAL S546 : STD_LOGIC;
    SIGNAL S547 : STD_LOGIC;
    SIGNAL S548 : STD_LOGIC;
    SIGNAL S549 : STD_LOGIC;
    SIGNAL S550 : STD_LOGIC;
    SIGNAL S551 : STD_LOGIC;
    SIGNAL S552 : STD_LOGIC;
    SIGNAL S553 : STD_LOGIC;
    SIGNAL S554 : STD_LOGIC;
    SIGNAL S555 : STD_LOGIC;
    SIGNAL S556 : STD_LOGIC;
    SIGNAL S557 : STD_LOGIC;
    SIGNAL S558 : STD_LOGIC;
    SIGNAL S559 : STD_LOGIC;
    SIGNAL S560 : STD_LOGIC;
    SIGNAL S561 : STD_LOGIC;
    SIGNAL S562 : STD_LOGIC;
    SIGNAL S563 : STD_LOGIC;
    SIGNAL S564 : STD_LOGIC;
    SIGNAL S565 : STD_LOGIC;
    SIGNAL S566 : STD_LOGIC;
    SIGNAL S567 : STD_LOGIC;
    SIGNAL S568 : STD_LOGIC;
    SIGNAL S569 : STD_LOGIC;
    SIGNAL S570 : STD_LOGIC;
    SIGNAL S571 : STD_LOGIC;
    SIGNAL S572 : STD_LOGIC;
    SIGNAL S573 : STD_LOGIC;
    SIGNAL S574 : STD_LOGIC;
    SIGNAL S575 : STD_LOGIC;
    SIGNAL S576 : STD_LOGIC;
    SIGNAL S577 : STD_LOGIC;
    SIGNAL S578 : STD_LOGIC;
    SIGNAL S579 : STD_LOGIC;
    SIGNAL S580 : STD_LOGIC;
    SIGNAL S581 : STD_LOGIC;
    SIGNAL S582 : STD_LOGIC;
    SIGNAL S583 : STD_LOGIC;
    SIGNAL S584 : STD_LOGIC;
    SIGNAL S585 : STD_LOGIC;
    SIGNAL S586 : STD_LOGIC;
    SIGNAL S587 : STD_LOGIC;
    SIGNAL S588 : STD_LOGIC;
    SIGNAL S589 : STD_LOGIC;
    SIGNAL S590 : STD_LOGIC;
    SIGNAL S591 : STD_LOGIC;
    SIGNAL S592 : STD_LOGIC;
    SIGNAL S593 : STD_LOGIC;
    SIGNAL S594 : STD_LOGIC;
    SIGNAL S595 : STD_LOGIC;
    SIGNAL S596 : STD_LOGIC;
    SIGNAL S597 : STD_LOGIC;
    SIGNAL S598 : STD_LOGIC;
    SIGNAL S599 : STD_LOGIC;
    SIGNAL S600 : STD_LOGIC;
    SIGNAL S601 : STD_LOGIC;
    SIGNAL S602 : STD_LOGIC;
    SIGNAL S603 : STD_LOGIC;
    SIGNAL S604 : STD_LOGIC;
    SIGNAL S605 : STD_LOGIC;
    SIGNAL S606 : STD_LOGIC;
    SIGNAL S607 : STD_LOGIC;
    SIGNAL S608 : STD_LOGIC;
    SIGNAL S609 : STD_LOGIC;
    SIGNAL S610 : STD_LOGIC;
    SIGNAL S611 : STD_LOGIC;
    SIGNAL S612 : STD_LOGIC;
    SIGNAL S613 : STD_LOGIC;
    SIGNAL S614 : STD_LOGIC;
    SIGNAL S615 : STD_LOGIC;
    SIGNAL S616 : STD_LOGIC;
    SIGNAL S617 : STD_LOGIC;
    SIGNAL S618 : STD_LOGIC;
    SIGNAL S619 : STD_LOGIC;
    SIGNAL S620 : STD_LOGIC;
    SIGNAL S621 : STD_LOGIC;
    SIGNAL S622 : STD_LOGIC;
    SIGNAL S623 : STD_LOGIC;
    SIGNAL S624 : STD_LOGIC;
    SIGNAL S625 : STD_LOGIC;
    SIGNAL S626 : STD_LOGIC;
    SIGNAL S627 : STD_LOGIC;
    SIGNAL S628 : STD_LOGIC;
    SIGNAL S629 : STD_LOGIC;
    SIGNAL S630 : STD_LOGIC;
    SIGNAL S631 : STD_LOGIC;
    SIGNAL S632 : STD_LOGIC;
    SIGNAL S633 : STD_LOGIC;
    SIGNAL S634 : STD_LOGIC;
    SIGNAL S635 : STD_LOGIC;
    SIGNAL S636 : STD_LOGIC;
    SIGNAL S637 : STD_LOGIC;
    SIGNAL S638 : STD_LOGIC;
    SIGNAL S639 : STD_LOGIC;
    SIGNAL S640 : STD_LOGIC;
    SIGNAL S641 : STD_LOGIC;
    SIGNAL S642 : STD_LOGIC;
    SIGNAL S643 : STD_LOGIC;
    SIGNAL S644 : STD_LOGIC;
    SIGNAL S645 : STD_LOGIC;
    SIGNAL S646 : STD_LOGIC;
    SIGNAL S647 : STD_LOGIC;
    SIGNAL S648 : STD_LOGIC;
    SIGNAL S649 : STD_LOGIC;
    SIGNAL S650 : STD_LOGIC;
    SIGNAL S651 : STD_LOGIC;
    SIGNAL S652 : STD_LOGIC;
    SIGNAL S653 : STD_LOGIC;
    SIGNAL S654 : STD_LOGIC;
    SIGNAL S655 : STD_LOGIC;
    SIGNAL S656 : STD_LOGIC;
    SIGNAL S657 : STD_LOGIC;
    SIGNAL S658 : STD_LOGIC;
    SIGNAL S659 : STD_LOGIC;
    SIGNAL S660 : STD_LOGIC;
    SIGNAL S661 : STD_LOGIC;
    SIGNAL S662 : STD_LOGIC;
    SIGNAL S663 : STD_LOGIC;
    SIGNAL S664 : STD_LOGIC;
    SIGNAL S665 : STD_LOGIC;
    SIGNAL S666 : STD_LOGIC;
    SIGNAL S667 : STD_LOGIC;
    SIGNAL S668 : STD_LOGIC;
    SIGNAL S669 : STD_LOGIC;
    SIGNAL S670 : STD_LOGIC;
    SIGNAL S671 : STD_LOGIC;
    SIGNAL S672 : STD_LOGIC;
    SIGNAL S673 : STD_LOGIC;
    SIGNAL S674 : STD_LOGIC;
    SIGNAL S675 : STD_LOGIC;
    SIGNAL S676 : STD_LOGIC;
    SIGNAL S677 : STD_LOGIC;
    SIGNAL S678 : STD_LOGIC;
    SIGNAL S679 : STD_LOGIC;
    SIGNAL S680 : STD_LOGIC;
    SIGNAL S681 : STD_LOGIC;
    SIGNAL S682 : STD_LOGIC;
    SIGNAL S683 : STD_LOGIC;
    SIGNAL S684 : STD_LOGIC;
    SIGNAL S685 : STD_LOGIC;
    SIGNAL S686 : STD_LOGIC;
    SIGNAL S687 : STD_LOGIC;
    SIGNAL S688 : STD_LOGIC;
    SIGNAL S689 : STD_LOGIC;
    SIGNAL S690 : STD_LOGIC;
    SIGNAL S691 : STD_LOGIC;
    SIGNAL S692 : STD_LOGIC;
    SIGNAL S693 : STD_LOGIC;
    SIGNAL S694 : STD_LOGIC;
    SIGNAL S695 : STD_LOGIC;
    SIGNAL S696 : STD_LOGIC;
    SIGNAL S697 : STD_LOGIC;
    SIGNAL S698 : STD_LOGIC;
    SIGNAL S699 : STD_LOGIC;
    SIGNAL S700 : STD_LOGIC;
    SIGNAL S701 : STD_LOGIC;
    SIGNAL S702 : STD_LOGIC;
    SIGNAL S703 : STD_LOGIC;
    SIGNAL S704 : STD_LOGIC;
    SIGNAL S705 : STD_LOGIC;
    SIGNAL S706 : STD_LOGIC;
    SIGNAL S707 : STD_LOGIC;
    SIGNAL S708 : STD_LOGIC;
    SIGNAL S709 : STD_LOGIC;
    SIGNAL S710 : STD_LOGIC;
    SIGNAL S711 : STD_LOGIC;
    SIGNAL S712 : STD_LOGIC;
    SIGNAL S713 : STD_LOGIC;
    SIGNAL S714 : STD_LOGIC;
    SIGNAL S715 : STD_LOGIC;
    SIGNAL S716 : STD_LOGIC;
    SIGNAL S717 : STD_LOGIC;
    SIGNAL S718 : STD_LOGIC;
    SIGNAL S719 : STD_LOGIC;
    SIGNAL S720 : STD_LOGIC;
    SIGNAL S721 : STD_LOGIC;
    SIGNAL S722 : STD_LOGIC;
    SIGNAL S723 : STD_LOGIC;
    SIGNAL S724 : STD_LOGIC;
    SIGNAL S725 : STD_LOGIC;
    SIGNAL S726 : STD_LOGIC;
    SIGNAL S727 : STD_LOGIC;
    SIGNAL S728 : STD_LOGIC;
    SIGNAL S729 : STD_LOGIC;
    SIGNAL S730 : STD_LOGIC;
    SIGNAL S731 : STD_LOGIC;
    SIGNAL S732 : STD_LOGIC;
    SIGNAL S733 : STD_LOGIC;
    SIGNAL S734 : STD_LOGIC;
    SIGNAL S735 : STD_LOGIC;
    SIGNAL S736 : STD_LOGIC;
    SIGNAL S737 : STD_LOGIC;
    SIGNAL S738 : STD_LOGIC;
    SIGNAL S739 : STD_LOGIC;
    SIGNAL S740 : STD_LOGIC;
    SIGNAL S741 : STD_LOGIC;
    SIGNAL S742 : STD_LOGIC;
    SIGNAL S743 : STD_LOGIC;
    SIGNAL S744 : STD_LOGIC;
    SIGNAL S745 : STD_LOGIC;
    SIGNAL S746 : STD_LOGIC;
    SIGNAL S747 : STD_LOGIC;
    SIGNAL S748 : STD_LOGIC;
    SIGNAL S749 : STD_LOGIC;
    SIGNAL S750 : STD_LOGIC;
    SIGNAL S751 : STD_LOGIC;
    SIGNAL S752 : STD_LOGIC;
    SIGNAL S753 : STD_LOGIC;
    SIGNAL S754 : STD_LOGIC;
    SIGNAL S755 : STD_LOGIC;
    SIGNAL S756 : STD_LOGIC;
    SIGNAL S757 : STD_LOGIC;
    SIGNAL S758 : STD_LOGIC;
    SIGNAL S759 : STD_LOGIC;
    SIGNAL S760 : STD_LOGIC;
    SIGNAL S761 : STD_LOGIC;
    SIGNAL S762 : STD_LOGIC;
    SIGNAL S763 : STD_LOGIC;
    SIGNAL S764 : STD_LOGIC;
    SIGNAL S765 : STD_LOGIC;
    SIGNAL S766 : STD_LOGIC;
    SIGNAL S767 : STD_LOGIC;
    SIGNAL S768 : STD_LOGIC;
    SIGNAL S769 : STD_LOGIC;
    SIGNAL S770 : STD_LOGIC;
    SIGNAL S771 : STD_LOGIC;
    SIGNAL S772 : STD_LOGIC;
    SIGNAL S773 : STD_LOGIC;
    SIGNAL S774 : STD_LOGIC;
    SIGNAL S775 : STD_LOGIC;
    SIGNAL S776 : STD_LOGIC;
    SIGNAL S777 : STD_LOGIC;
    SIGNAL S778 : STD_LOGIC;
    SIGNAL S779 : STD_LOGIC;
    SIGNAL S780 : STD_LOGIC;
    SIGNAL S781 : STD_LOGIC;
    SIGNAL S782 : STD_LOGIC;
    SIGNAL S783 : STD_LOGIC;
    SIGNAL S784 : STD_LOGIC;
    SIGNAL S785 : STD_LOGIC;
    SIGNAL S786 : STD_LOGIC;
    SIGNAL S787 : STD_LOGIC;
    SIGNAL S788 : STD_LOGIC;
    SIGNAL S789 : STD_LOGIC;
    SIGNAL S790 : STD_LOGIC;
    SIGNAL S791 : STD_LOGIC;
    SIGNAL S792 : STD_LOGIC;
    SIGNAL S793 : STD_LOGIC;
    SIGNAL S794 : STD_LOGIC;
    SIGNAL S795 : STD_LOGIC;
    SIGNAL S796 : STD_LOGIC;
    SIGNAL S797 : STD_LOGIC;
    SIGNAL S798 : STD_LOGIC;
    SIGNAL S799 : STD_LOGIC;
    SIGNAL S800 : STD_LOGIC;
    SIGNAL S801 : STD_LOGIC;
    SIGNAL S802 : STD_LOGIC;
    SIGNAL S803 : STD_LOGIC;
    SIGNAL S804 : STD_LOGIC;
    SIGNAL S805 : STD_LOGIC;
    SIGNAL S806 : STD_LOGIC;
    SIGNAL S807 : STD_LOGIC;
    SIGNAL S808 : STD_LOGIC;
    SIGNAL S809 : STD_LOGIC;
    SIGNAL S810 : STD_LOGIC;
    SIGNAL S811 : STD_LOGIC;
    SIGNAL S812 : STD_LOGIC;
    SIGNAL S813 : STD_LOGIC;
    SIGNAL S814 : STD_LOGIC;
    SIGNAL S815 : STD_LOGIC;
    SIGNAL S816 : STD_LOGIC;
    SIGNAL S817 : STD_LOGIC;
    SIGNAL S818 : STD_LOGIC;
    SIGNAL S819 : STD_LOGIC;
    SIGNAL S820 : STD_LOGIC;
    SIGNAL S821 : STD_LOGIC;
    SIGNAL S822 : STD_LOGIC;
    SIGNAL S823 : STD_LOGIC;
    SIGNAL S824 : STD_LOGIC;
    SIGNAL S825 : STD_LOGIC;
    SIGNAL S826 : STD_LOGIC;
    SIGNAL S827 : STD_LOGIC;
    SIGNAL S828 : STD_LOGIC;
    SIGNAL S829 : STD_LOGIC;
    SIGNAL S830 : STD_LOGIC;
    SIGNAL S831 : STD_LOGIC;
    SIGNAL S832 : STD_LOGIC;
    SIGNAL S833 : STD_LOGIC;
    SIGNAL S834 : STD_LOGIC;
    SIGNAL S835 : STD_LOGIC;
    SIGNAL S836 : STD_LOGIC;
    SIGNAL S837 : STD_LOGIC;
    SIGNAL S838 : STD_LOGIC;
    SIGNAL S839 : STD_LOGIC;
    SIGNAL S840 : STD_LOGIC;
    SIGNAL S841 : STD_LOGIC;
    SIGNAL S842 : STD_LOGIC;
    SIGNAL S843 : STD_LOGIC;
    SIGNAL S844 : STD_LOGIC;
    SIGNAL S845 : STD_LOGIC;
    SIGNAL S846 : STD_LOGIC;
    SIGNAL S847 : STD_LOGIC;
    SIGNAL S848 : STD_LOGIC;
    SIGNAL S849 : STD_LOGIC;
    SIGNAL S850 : STD_LOGIC;
    SIGNAL S851 : STD_LOGIC;
    SIGNAL S852 : STD_LOGIC;
    SIGNAL S853 : STD_LOGIC;
    SIGNAL S854 : STD_LOGIC;
    SIGNAL S855 : STD_LOGIC;
    SIGNAL S856 : STD_LOGIC;
    SIGNAL S857 : STD_LOGIC;
    SIGNAL S858 : STD_LOGIC;
    SIGNAL S859 : STD_LOGIC;
    SIGNAL S860 : STD_LOGIC;
    SIGNAL S861 : STD_LOGIC;
    SIGNAL S862 : STD_LOGIC;
    SIGNAL S863 : STD_LOGIC;
    SIGNAL S864 : STD_LOGIC;
    SIGNAL S865 : STD_LOGIC;
    SIGNAL S866 : STD_LOGIC;
    SIGNAL S867 : STD_LOGIC;
    SIGNAL S868 : STD_LOGIC;
    SIGNAL S869 : STD_LOGIC;
    SIGNAL S870 : STD_LOGIC;
    SIGNAL S871 : STD_LOGIC;
    SIGNAL S872 : STD_LOGIC;
    SIGNAL S873 : STD_LOGIC;
    SIGNAL S874 : STD_LOGIC;
    SIGNAL S875 : STD_LOGIC;
    SIGNAL S876 : STD_LOGIC;
    SIGNAL S877 : STD_LOGIC;
    SIGNAL S878 : STD_LOGIC;
    SIGNAL S879 : STD_LOGIC;
    SIGNAL S880 : STD_LOGIC;
    SIGNAL S881 : STD_LOGIC;
    SIGNAL S882 : STD_LOGIC;
    SIGNAL S883 : STD_LOGIC;
    SIGNAL S884 : STD_LOGIC;
    SIGNAL S885 : STD_LOGIC;
    SIGNAL S886 : STD_LOGIC;
    SIGNAL S887 : STD_LOGIC;
    SIGNAL S888 : STD_LOGIC;
    SIGNAL S889 : STD_LOGIC;
    SIGNAL S890 : STD_LOGIC;
    SIGNAL S891 : STD_LOGIC;
    SIGNAL S892 : STD_LOGIC;
    SIGNAL S893 : STD_LOGIC;
    SIGNAL S894 : STD_LOGIC;
    SIGNAL S895 : STD_LOGIC;
    SIGNAL S896 : STD_LOGIC;
    SIGNAL S897 : STD_LOGIC;
    SIGNAL S898 : STD_LOGIC;
    SIGNAL S899 : STD_LOGIC;
    SIGNAL S900 : STD_LOGIC;
    SIGNAL S901 : STD_LOGIC;
    SIGNAL S902 : STD_LOGIC;
    SIGNAL S903 : STD_LOGIC;
    SIGNAL S904 : STD_LOGIC;
    SIGNAL S905 : STD_LOGIC;
    SIGNAL S906 : STD_LOGIC;
    SIGNAL S907 : STD_LOGIC;
    SIGNAL S908 : STD_LOGIC;
    SIGNAL S909 : STD_LOGIC;
    SIGNAL S910 : STD_LOGIC;
    SIGNAL S911 : STD_LOGIC;
    SIGNAL S912 : STD_LOGIC;
    SIGNAL S913 : STD_LOGIC;
    SIGNAL S914 : STD_LOGIC;
    SIGNAL S915 : STD_LOGIC;
    SIGNAL S916 : STD_LOGIC;
    SIGNAL S917 : STD_LOGIC;
    SIGNAL S918 : STD_LOGIC;
    SIGNAL S919 : STD_LOGIC;
    SIGNAL S920 : STD_LOGIC;
    SIGNAL S921 : STD_LOGIC;
    SIGNAL S922 : STD_LOGIC;
    SIGNAL S923 : STD_LOGIC;
    SIGNAL S924 : STD_LOGIC;
    SIGNAL S925 : STD_LOGIC;
    SIGNAL S926 : STD_LOGIC;
    SIGNAL S927 : STD_LOGIC;
    SIGNAL S928 : STD_LOGIC;
    SIGNAL S929 : STD_LOGIC;
    SIGNAL S930 : STD_LOGIC;
    SIGNAL S931 : STD_LOGIC;
    SIGNAL S932 : STD_LOGIC;
    SIGNAL S933 : STD_LOGIC;
    SIGNAL S934 : STD_LOGIC;
    SIGNAL S935 : STD_LOGIC;
    SIGNAL S936 : STD_LOGIC;
    SIGNAL S937 : STD_LOGIC;
    SIGNAL S938 : STD_LOGIC;
    SIGNAL S939 : STD_LOGIC;
    SIGNAL S940 : STD_LOGIC;
    SIGNAL S941 : STD_LOGIC;
    SIGNAL S942 : STD_LOGIC;
    SIGNAL S943 : STD_LOGIC;
    SIGNAL S944 : STD_LOGIC;
    SIGNAL S945 : STD_LOGIC;
    SIGNAL S946 : STD_LOGIC;
    SIGNAL S947 : STD_LOGIC;
    SIGNAL S948 : STD_LOGIC;
    SIGNAL S949 : STD_LOGIC;
    SIGNAL S950 : STD_LOGIC;
    SIGNAL S951 : STD_LOGIC;
    SIGNAL S952 : STD_LOGIC;
    SIGNAL S953 : STD_LOGIC;
    SIGNAL S954 : STD_LOGIC;
    SIGNAL S955 : STD_LOGIC;
    SIGNAL S956 : STD_LOGIC;
    SIGNAL S957 : STD_LOGIC;
    SIGNAL S958 : STD_LOGIC;
    SIGNAL S959 : STD_LOGIC;
    SIGNAL S960 : STD_LOGIC;
    SIGNAL S961 : STD_LOGIC;
    SIGNAL S962 : STD_LOGIC;
    SIGNAL S963 : STD_LOGIC;
    SIGNAL S964 : STD_LOGIC;
    SIGNAL S965 : STD_LOGIC;
    SIGNAL S966 : STD_LOGIC;
    SIGNAL S967 : STD_LOGIC;
    SIGNAL S968 : STD_LOGIC;
    SIGNAL S969 : STD_LOGIC;
    SIGNAL S970 : STD_LOGIC;
    SIGNAL S971 : STD_LOGIC;
    SIGNAL S972 : STD_LOGIC;
    SIGNAL S973 : STD_LOGIC;
    SIGNAL S974 : STD_LOGIC;
    SIGNAL S975 : STD_LOGIC;
    SIGNAL S976 : STD_LOGIC;
    SIGNAL S977 : STD_LOGIC;
    SIGNAL S978 : STD_LOGIC;
    SIGNAL S979 : STD_LOGIC;
    SIGNAL S980 : STD_LOGIC;
    SIGNAL S981 : STD_LOGIC;
    SIGNAL S982 : STD_LOGIC;
    SIGNAL S983 : STD_LOGIC;
    SIGNAL S984 : STD_LOGIC;
    SIGNAL S985 : STD_LOGIC;
    SIGNAL S986 : STD_LOGIC;
    SIGNAL S987 : STD_LOGIC;
    SIGNAL S988 : STD_LOGIC;
    SIGNAL S989 : STD_LOGIC;
    SIGNAL S990 : STD_LOGIC;
    SIGNAL S991 : STD_LOGIC;
    SIGNAL S992 : STD_LOGIC;
    SIGNAL S993 : STD_LOGIC;
    SIGNAL S994 : STD_LOGIC;
    SIGNAL S995 : STD_LOGIC;
    SIGNAL S996 : STD_LOGIC;
    SIGNAL S997 : STD_LOGIC;
    SIGNAL S998 : STD_LOGIC;
    SIGNAL S999 : STD_LOGIC;
    SIGNAL S1000 : STD_LOGIC;
    SIGNAL S1001 : STD_LOGIC;
    SIGNAL S1002 : STD_LOGIC;
    SIGNAL S1003 : STD_LOGIC;
    SIGNAL S1004 : STD_LOGIC;
    SIGNAL S1005 : STD_LOGIC;
    SIGNAL S1006 : STD_LOGIC;
    SIGNAL S1007 : STD_LOGIC;
    SIGNAL S1008 : STD_LOGIC;
    SIGNAL S1009 : STD_LOGIC;
    SIGNAL S1010 : STD_LOGIC;
    SIGNAL S1011 : STD_LOGIC;
    SIGNAL S1012 : STD_LOGIC;
    SIGNAL S1013 : STD_LOGIC;
    SIGNAL S1014 : STD_LOGIC;
    SIGNAL S1015 : STD_LOGIC;
    SIGNAL S1016 : STD_LOGIC;
    SIGNAL S1017 : STD_LOGIC;
    SIGNAL S1018 : STD_LOGIC;
    SIGNAL S1019 : STD_LOGIC;
    SIGNAL S1020 : STD_LOGIC;
    SIGNAL S1021 : STD_LOGIC;
    SIGNAL S1022 : STD_LOGIC;
    SIGNAL S1023 : STD_LOGIC;
    SIGNAL S1024 : STD_LOGIC;
    SIGNAL S1025 : STD_LOGIC;
    SIGNAL S1026 : STD_LOGIC;
    SIGNAL S1027 : STD_LOGIC;
    SIGNAL S1028 : STD_LOGIC;
    SIGNAL S1029 : STD_LOGIC;
    SIGNAL S1030 : STD_LOGIC;
    SIGNAL S1031 : STD_LOGIC;
    SIGNAL S1032 : STD_LOGIC;
    SIGNAL S1033 : STD_LOGIC;
    SIGNAL S1034 : STD_LOGIC;
    SIGNAL S1035 : STD_LOGIC;
    SIGNAL S1036 : STD_LOGIC;
    SIGNAL S1037 : STD_LOGIC;
    SIGNAL S1038 : STD_LOGIC;
    SIGNAL S1039 : STD_LOGIC;
    SIGNAL S1040 : STD_LOGIC;
    SIGNAL S1041 : STD_LOGIC;
    SIGNAL S1042 : STD_LOGIC;
    SIGNAL S1043 : STD_LOGIC;
    SIGNAL S1044 : STD_LOGIC;
    SIGNAL S1045 : STD_LOGIC;
    SIGNAL S1046 : STD_LOGIC;
    SIGNAL S1047 : STD_LOGIC;
    SIGNAL S1048 : STD_LOGIC;
    SIGNAL S1049 : STD_LOGIC;
    SIGNAL S1050 : STD_LOGIC;
    SIGNAL S1051 : STD_LOGIC;
    SIGNAL S1052 : STD_LOGIC;
    SIGNAL S1053 : STD_LOGIC;
    SIGNAL S1054 : STD_LOGIC;
    SIGNAL S1055 : STD_LOGIC;
    SIGNAL S1056 : STD_LOGIC;
    SIGNAL S1057 : STD_LOGIC;
    SIGNAL S1058 : STD_LOGIC;
    SIGNAL S1059 : STD_LOGIC;
    SIGNAL S1060 : STD_LOGIC;
    SIGNAL S1061 : STD_LOGIC;
    SIGNAL S1062 : STD_LOGIC;
    SIGNAL S1063 : STD_LOGIC;
    SIGNAL S1064 : STD_LOGIC;
    SIGNAL S1065 : STD_LOGIC;
    SIGNAL S1066 : STD_LOGIC;
    SIGNAL S1067 : STD_LOGIC;
    SIGNAL S1068 : STD_LOGIC;
    SIGNAL S1069 : STD_LOGIC;
    SIGNAL S1070 : STD_LOGIC;
    SIGNAL S1071 : STD_LOGIC;
    SIGNAL S1072 : STD_LOGIC;
    SIGNAL S1073 : STD_LOGIC;
    SIGNAL S1074 : STD_LOGIC;
    SIGNAL S1075 : STD_LOGIC;
    SIGNAL S1076 : STD_LOGIC;
    SIGNAL S1077 : STD_LOGIC;
    SIGNAL S1078 : STD_LOGIC;
    SIGNAL S1079 : STD_LOGIC;
    SIGNAL S1080 : STD_LOGIC;
    SIGNAL S1081 : STD_LOGIC;
    SIGNAL S1082 : STD_LOGIC;
    SIGNAL S1083 : STD_LOGIC;
    SIGNAL S1084 : STD_LOGIC;
    SIGNAL S1085 : STD_LOGIC;
    SIGNAL S1086 : STD_LOGIC;
    SIGNAL S1087 : STD_LOGIC;
    SIGNAL S1088 : STD_LOGIC;
    SIGNAL S1089 : STD_LOGIC;
    SIGNAL S1090 : STD_LOGIC;
    SIGNAL S1091 : STD_LOGIC;
    SIGNAL S1092 : STD_LOGIC;
    SIGNAL S1093 : STD_LOGIC;
    SIGNAL S1094 : STD_LOGIC;
    SIGNAL S1095 : STD_LOGIC;
    SIGNAL S1096 : STD_LOGIC;
    SIGNAL S1097 : STD_LOGIC;
    SIGNAL S1098 : STD_LOGIC;
    SIGNAL S1099 : STD_LOGIC;
    SIGNAL S1100 : STD_LOGIC;
    SIGNAL S1101 : STD_LOGIC;
    SIGNAL S1102 : STD_LOGIC;
    SIGNAL S1103 : STD_LOGIC;
    SIGNAL S1104 : STD_LOGIC;
    SIGNAL S1105 : STD_LOGIC;
    SIGNAL S1106 : STD_LOGIC;
    SIGNAL S1107 : STD_LOGIC;
    SIGNAL S1108 : STD_LOGIC;
    SIGNAL S1109 : STD_LOGIC;
    SIGNAL S1110 : STD_LOGIC;
    SIGNAL S1111 : STD_LOGIC;
    SIGNAL S1112 : STD_LOGIC;
    SIGNAL S1113 : STD_LOGIC;
    SIGNAL S1114 : STD_LOGIC;
    SIGNAL S1115 : STD_LOGIC;
    SIGNAL S1116 : STD_LOGIC;
    SIGNAL S1117 : STD_LOGIC;
    SIGNAL S1118 : STD_LOGIC;
    SIGNAL S1119 : STD_LOGIC;
    SIGNAL S1120 : STD_LOGIC;
    SIGNAL S1121 : STD_LOGIC;
    SIGNAL S1122 : STD_LOGIC;
    SIGNAL S1123 : STD_LOGIC;
    SIGNAL S1124 : STD_LOGIC;
    SIGNAL S1125 : STD_LOGIC;
    SIGNAL S1126 : STD_LOGIC;
    SIGNAL S1127 : STD_LOGIC;
    SIGNAL S1128 : STD_LOGIC;
    SIGNAL S1129 : STD_LOGIC;
    SIGNAL S1130 : STD_LOGIC;
    SIGNAL S1131 : STD_LOGIC;
    SIGNAL S1132 : STD_LOGIC;
    SIGNAL S1133 : STD_LOGIC;
    SIGNAL S1134 : STD_LOGIC;
    SIGNAL S1135 : STD_LOGIC;
    SIGNAL S1136 : STD_LOGIC;
    SIGNAL S1137 : STD_LOGIC;
    SIGNAL S1138 : STD_LOGIC;
    SIGNAL S1139 : STD_LOGIC;
    SIGNAL S1140 : STD_LOGIC;
    SIGNAL S1141 : STD_LOGIC;
    SIGNAL S1142 : STD_LOGIC;
    SIGNAL S1143 : STD_LOGIC;
    SIGNAL S1144 : STD_LOGIC;
    SIGNAL S1145 : STD_LOGIC;
    SIGNAL S1146 : STD_LOGIC;
    SIGNAL S1147 : STD_LOGIC;
    SIGNAL S1148 : STD_LOGIC;
    SIGNAL S1149 : STD_LOGIC;
    SIGNAL S1150 : STD_LOGIC;
    SIGNAL S1151 : STD_LOGIC;
    SIGNAL S1152 : STD_LOGIC;
    SIGNAL S1153 : STD_LOGIC;
    SIGNAL S1154 : STD_LOGIC;
    SIGNAL S1155 : STD_LOGIC;
    SIGNAL S1156 : STD_LOGIC;
    SIGNAL S1157 : STD_LOGIC;
    SIGNAL S1158 : STD_LOGIC;
    SIGNAL S1159 : STD_LOGIC;
    SIGNAL S1160 : STD_LOGIC;
    SIGNAL S1161 : STD_LOGIC;
    SIGNAL S1162 : STD_LOGIC;
    SIGNAL S1163 : STD_LOGIC;
    SIGNAL S1164 : STD_LOGIC;
    SIGNAL S1165 : STD_LOGIC;
    SIGNAL S1166 : STD_LOGIC;
    SIGNAL S1167 : STD_LOGIC;
    SIGNAL S1168 : STD_LOGIC;
    SIGNAL S1169 : STD_LOGIC;
    SIGNAL S1170 : STD_LOGIC;
    SIGNAL S1171 : STD_LOGIC;
    SIGNAL S1172 : STD_LOGIC;
    SIGNAL S1173 : STD_LOGIC;
    SIGNAL S1174 : STD_LOGIC;
    SIGNAL S1175 : STD_LOGIC;
    SIGNAL S1176 : STD_LOGIC;
    SIGNAL S1177 : STD_LOGIC;
    SIGNAL S1178 : STD_LOGIC;
    SIGNAL S1179 : STD_LOGIC;
    SIGNAL S1180 : STD_LOGIC;
    SIGNAL S1181 : STD_LOGIC;
    SIGNAL S1182 : STD_LOGIC;
    SIGNAL S1183 : STD_LOGIC;
    SIGNAL S1184 : STD_LOGIC;
    SIGNAL S1185 : STD_LOGIC;
    SIGNAL S1186 : STD_LOGIC;
    SIGNAL S1187 : STD_LOGIC;
    SIGNAL S1188 : STD_LOGIC;
    SIGNAL S1189 : STD_LOGIC;
    SIGNAL S1190 : STD_LOGIC;
    SIGNAL S1191 : STD_LOGIC;
    SIGNAL S1192 : STD_LOGIC;
    SIGNAL S1193 : STD_LOGIC;
    SIGNAL S1194 : STD_LOGIC;
    SIGNAL S1195 : STD_LOGIC;
    SIGNAL S1196 : STD_LOGIC;
    SIGNAL S1197 : STD_LOGIC;
    SIGNAL S1198 : STD_LOGIC;
    SIGNAL S1199 : STD_LOGIC;
    SIGNAL S1200 : STD_LOGIC;
    SIGNAL S1201 : STD_LOGIC;
    SIGNAL S1202 : STD_LOGIC;
    SIGNAL S1203 : STD_LOGIC;
    SIGNAL S1204 : STD_LOGIC;
    SIGNAL S1205 : STD_LOGIC;
    SIGNAL S1206 : STD_LOGIC;
    SIGNAL S1207 : STD_LOGIC;
    SIGNAL S1208 : STD_LOGIC;
    SIGNAL S1209 : STD_LOGIC;
    SIGNAL S1210 : STD_LOGIC;
    SIGNAL S1211 : STD_LOGIC;
    SIGNAL S1212 : STD_LOGIC;
    SIGNAL S1213 : STD_LOGIC;
    SIGNAL S1214 : STD_LOGIC;
    SIGNAL S1215 : STD_LOGIC;
    SIGNAL S1216 : STD_LOGIC;
    SIGNAL S1217 : STD_LOGIC;
    SIGNAL S1218 : STD_LOGIC;
    SIGNAL S1219 : STD_LOGIC;
    SIGNAL S1220 : STD_LOGIC;
    SIGNAL S1221 : STD_LOGIC;
    SIGNAL S1222 : STD_LOGIC;
    SIGNAL S1223 : STD_LOGIC;
    SIGNAL S1224 : STD_LOGIC;
    SIGNAL S1225 : STD_LOGIC;
    SIGNAL S1226 : STD_LOGIC;
    SIGNAL S1227 : STD_LOGIC;
    SIGNAL S1228 : STD_LOGIC;
    SIGNAL S1229 : STD_LOGIC;
    SIGNAL S1230 : STD_LOGIC;
    SIGNAL S1231 : STD_LOGIC;
    SIGNAL S1232 : STD_LOGIC;
    SIGNAL S1233 : STD_LOGIC;
    SIGNAL S1234 : STD_LOGIC;
    SIGNAL S1235 : STD_LOGIC;
    SIGNAL S1236 : STD_LOGIC;
    SIGNAL S1237 : STD_LOGIC;
    SIGNAL S1238 : STD_LOGIC;
    SIGNAL S1239 : STD_LOGIC;
    SIGNAL S1240 : STD_LOGIC;
    SIGNAL S1241 : STD_LOGIC;
    SIGNAL S1242 : STD_LOGIC;
    SIGNAL S1243 : STD_LOGIC;
    SIGNAL S1244 : STD_LOGIC;
    SIGNAL S1245 : STD_LOGIC;
    SIGNAL S1246 : STD_LOGIC;
    SIGNAL S1247 : STD_LOGIC;
    SIGNAL S1248 : STD_LOGIC;
    SIGNAL S1249 : STD_LOGIC;
    SIGNAL S1250 : STD_LOGIC;
    SIGNAL S1251 : STD_LOGIC;
    SIGNAL S1252 : STD_LOGIC;
    SIGNAL S1253 : STD_LOGIC;
    SIGNAL S1254 : STD_LOGIC;
    SIGNAL S1255 : STD_LOGIC;
    SIGNAL S1256 : STD_LOGIC;
    SIGNAL S1257 : STD_LOGIC;
    SIGNAL S1258 : STD_LOGIC;
    SIGNAL S1259 : STD_LOGIC;
    SIGNAL S1260 : STD_LOGIC;
    SIGNAL S1261 : STD_LOGIC;
    SIGNAL S1262 : STD_LOGIC;
    SIGNAL S1263 : STD_LOGIC;
    SIGNAL S1264 : STD_LOGIC;
    SIGNAL S1265 : STD_LOGIC;
    SIGNAL S1266 : STD_LOGIC;
    SIGNAL S1267 : STD_LOGIC;
    SIGNAL S1268 : STD_LOGIC;
    SIGNAL S1269 : STD_LOGIC;
    SIGNAL S1270 : STD_LOGIC;
    SIGNAL S1271 : STD_LOGIC;
    SIGNAL S1272 : STD_LOGIC;
    SIGNAL S1273 : STD_LOGIC;
    SIGNAL S1274 : STD_LOGIC;
    SIGNAL S1275 : STD_LOGIC;
    SIGNAL S1276 : STD_LOGIC;
    SIGNAL S1277 : STD_LOGIC;
    SIGNAL S1278 : STD_LOGIC;
    SIGNAL S1279 : STD_LOGIC;
    SIGNAL S1280 : STD_LOGIC;
    SIGNAL S1281 : STD_LOGIC;
    SIGNAL S1282 : STD_LOGIC;
    SIGNAL S1283 : STD_LOGIC;
    SIGNAL S1284 : STD_LOGIC;
    SIGNAL S1285 : STD_LOGIC;
    SIGNAL S1286 : STD_LOGIC;
    SIGNAL S1287 : STD_LOGIC;
    SIGNAL S1288 : STD_LOGIC;
    SIGNAL S1289 : STD_LOGIC;
    SIGNAL S1290 : STD_LOGIC;
    SIGNAL S1291 : STD_LOGIC;
    SIGNAL S1292 : STD_LOGIC;
    SIGNAL S1293 : STD_LOGIC;
    SIGNAL S1294 : STD_LOGIC;
    SIGNAL S1295 : STD_LOGIC;
    SIGNAL S1296 : STD_LOGIC;
    SIGNAL S1297 : STD_LOGIC;
    SIGNAL S1298 : STD_LOGIC;
    SIGNAL S1299 : STD_LOGIC;
    SIGNAL S1300 : STD_LOGIC;
    SIGNAL S1301 : STD_LOGIC;
    SIGNAL S1302 : STD_LOGIC;
    SIGNAL S1303 : STD_LOGIC;
    SIGNAL S1304 : STD_LOGIC;
    SIGNAL S1305 : STD_LOGIC;
    SIGNAL S1306 : STD_LOGIC;
    SIGNAL S1307 : STD_LOGIC;
    SIGNAL S1308 : STD_LOGIC;
    SIGNAL S1309 : STD_LOGIC;
    SIGNAL S1310 : STD_LOGIC;
    SIGNAL S1311 : STD_LOGIC;
    SIGNAL S1312 : STD_LOGIC;
    SIGNAL S1313 : STD_LOGIC;
    SIGNAL S1314 : STD_LOGIC;
    SIGNAL S1315 : STD_LOGIC;
    SIGNAL S1316 : STD_LOGIC;
    SIGNAL S1317 : STD_LOGIC;
    SIGNAL S1318 : STD_LOGIC;
    SIGNAL S1319 : STD_LOGIC;
    SIGNAL S1320 : STD_LOGIC;
    SIGNAL S1321 : STD_LOGIC;
    SIGNAL S1322 : STD_LOGIC;
    SIGNAL S1323 : STD_LOGIC;
    SIGNAL S1324 : STD_LOGIC;
    SIGNAL S1325 : STD_LOGIC;
    SIGNAL S1326 : STD_LOGIC;
    SIGNAL S1327 : STD_LOGIC;
    SIGNAL S1328 : STD_LOGIC;
    SIGNAL S1329 : STD_LOGIC;
    SIGNAL S1330 : STD_LOGIC;
    SIGNAL S1331 : STD_LOGIC;
    SIGNAL S1332 : STD_LOGIC;
    SIGNAL S1333 : STD_LOGIC;
    SIGNAL S1334 : STD_LOGIC;
    SIGNAL S1335 : STD_LOGIC;
    SIGNAL S1336 : STD_LOGIC;
    SIGNAL S1337 : STD_LOGIC;
    SIGNAL S1338 : STD_LOGIC;
    SIGNAL S1339 : STD_LOGIC;
    SIGNAL S1340 : STD_LOGIC;
    SIGNAL S1341 : STD_LOGIC;
    SIGNAL S1342 : STD_LOGIC;
    SIGNAL S1343 : STD_LOGIC;
    SIGNAL S1344 : STD_LOGIC;
    SIGNAL S1345 : STD_LOGIC;
    SIGNAL S1346 : STD_LOGIC;
    SIGNAL S1347 : STD_LOGIC;
    SIGNAL S1348 : STD_LOGIC;
    SIGNAL S1349 : STD_LOGIC;
    SIGNAL S1350 : STD_LOGIC;
    SIGNAL S1351 : STD_LOGIC;
    SIGNAL S1352 : STD_LOGIC;
    SIGNAL S1353 : STD_LOGIC;
    SIGNAL S1354 : STD_LOGIC;
    SIGNAL S1355 : STD_LOGIC;
    SIGNAL S1356 : STD_LOGIC;
    SIGNAL S1357 : STD_LOGIC;
    SIGNAL S1358 : STD_LOGIC;
    SIGNAL S1359 : STD_LOGIC;
    SIGNAL S1360 : STD_LOGIC;
    SIGNAL S1361 : STD_LOGIC;
    SIGNAL S1362 : STD_LOGIC;
    SIGNAL S1363 : STD_LOGIC;
    SIGNAL S1364 : STD_LOGIC;
    SIGNAL S1365 : STD_LOGIC;
    SIGNAL S1366 : STD_LOGIC;
    SIGNAL S1367 : STD_LOGIC;
    SIGNAL S1368 : STD_LOGIC;
    SIGNAL S1369 : STD_LOGIC;
    SIGNAL S1370 : STD_LOGIC;
    SIGNAL S1371 : STD_LOGIC;
    SIGNAL S1372 : STD_LOGIC;
    SIGNAL S1373 : STD_LOGIC;
    SIGNAL S1374 : STD_LOGIC;
    SIGNAL S1375 : STD_LOGIC;
    SIGNAL S1376 : STD_LOGIC;
    SIGNAL S1377 : STD_LOGIC;
    SIGNAL S1378 : STD_LOGIC;
    SIGNAL S1379 : STD_LOGIC;
    SIGNAL S1380 : STD_LOGIC;
    SIGNAL S1381 : STD_LOGIC;
    SIGNAL S1382 : STD_LOGIC;
    SIGNAL S1383 : STD_LOGIC;
    SIGNAL S1384 : STD_LOGIC;
    SIGNAL S1385 : STD_LOGIC;
    SIGNAL S1386 : STD_LOGIC;
    SIGNAL S1387 : STD_LOGIC;
    SIGNAL S1388 : STD_LOGIC;
    SIGNAL S1389 : STD_LOGIC;
    SIGNAL S1390 : STD_LOGIC;
    SIGNAL S1391 : STD_LOGIC;
    SIGNAL S1392 : STD_LOGIC;
    SIGNAL S1393 : STD_LOGIC;
    SIGNAL S1394 : STD_LOGIC;
    SIGNAL S1395 : STD_LOGIC;
    SIGNAL S1396 : STD_LOGIC;
    SIGNAL S1397 : STD_LOGIC;
    SIGNAL S1398 : STD_LOGIC;
    SIGNAL S1399 : STD_LOGIC;
    SIGNAL S1400 : STD_LOGIC;
    SIGNAL S1401 : STD_LOGIC;
    SIGNAL S1402 : STD_LOGIC;
    SIGNAL S1403 : STD_LOGIC;
    SIGNAL S1404 : STD_LOGIC;
    SIGNAL S1405 : STD_LOGIC;
    SIGNAL S1406 : STD_LOGIC;
    SIGNAL S1407 : STD_LOGIC;
    SIGNAL S1408 : STD_LOGIC;
    SIGNAL S1409 : STD_LOGIC;
    SIGNAL S1410 : STD_LOGIC;
    SIGNAL S1411 : STD_LOGIC;
    SIGNAL S1412 : STD_LOGIC;
    SIGNAL S1413 : STD_LOGIC;
    SIGNAL S1414 : STD_LOGIC;
    SIGNAL S1415 : STD_LOGIC;
    SIGNAL S1416 : STD_LOGIC;
    SIGNAL S1417 : STD_LOGIC;
    SIGNAL S1418 : STD_LOGIC;
    SIGNAL S1419 : STD_LOGIC;
    SIGNAL S1420 : STD_LOGIC;
    SIGNAL S1421 : STD_LOGIC;
    SIGNAL S1422 : STD_LOGIC;
    SIGNAL S1423 : STD_LOGIC;
    SIGNAL S1424 : STD_LOGIC;
    SIGNAL S1425 : STD_LOGIC;
    SIGNAL S1426 : STD_LOGIC;
    SIGNAL S1427 : STD_LOGIC;
    SIGNAL S1428 : STD_LOGIC;
    SIGNAL S1429 : STD_LOGIC;
    SIGNAL S1430 : STD_LOGIC;
    SIGNAL S1431 : STD_LOGIC;
    SIGNAL S1432 : STD_LOGIC;
    SIGNAL S1433 : STD_LOGIC;
    SIGNAL S1434 : STD_LOGIC;
    SIGNAL S1435 : STD_LOGIC;
    SIGNAL S1436 : STD_LOGIC;
    SIGNAL S1437 : STD_LOGIC;
    SIGNAL S1438 : STD_LOGIC;
    SIGNAL S1439 : STD_LOGIC;
    SIGNAL S1440 : STD_LOGIC;
    SIGNAL S1441 : STD_LOGIC;
    SIGNAL S1442 : STD_LOGIC;
    SIGNAL S1443 : STD_LOGIC;
    SIGNAL S1444 : STD_LOGIC;
    SIGNAL S1445 : STD_LOGIC;
    SIGNAL S1446 : STD_LOGIC;
    SIGNAL S1447 : STD_LOGIC;
    SIGNAL S1448 : STD_LOGIC;
    SIGNAL S1449 : STD_LOGIC;
    SIGNAL S1450 : STD_LOGIC;
    SIGNAL S1451 : STD_LOGIC;
    SIGNAL S1452 : STD_LOGIC;
    SIGNAL S1453 : STD_LOGIC;
    SIGNAL S1454 : STD_LOGIC;
    SIGNAL S1455 : STD_LOGIC;
    SIGNAL S1456 : STD_LOGIC;
    SIGNAL S1457 : STD_LOGIC;
    SIGNAL S1458 : STD_LOGIC;
    SIGNAL S1459 : STD_LOGIC;
    SIGNAL S1460 : STD_LOGIC;
    SIGNAL S1461 : STD_LOGIC;
    SIGNAL S1462 : STD_LOGIC;
    SIGNAL S1463 : STD_LOGIC;
    SIGNAL S1464 : STD_LOGIC;
    SIGNAL S1465 : STD_LOGIC;
    SIGNAL S1466 : STD_LOGIC;
    SIGNAL S1467 : STD_LOGIC;
    SIGNAL S1468 : STD_LOGIC;
    SIGNAL S1469 : STD_LOGIC;
    SIGNAL S1470 : STD_LOGIC;
    SIGNAL S1471 : STD_LOGIC;
    SIGNAL S1472 : STD_LOGIC;
    SIGNAL S1473 : STD_LOGIC;
    SIGNAL S1474 : STD_LOGIC;
    SIGNAL S1475 : STD_LOGIC;
    SIGNAL S1476 : STD_LOGIC;
    SIGNAL S1477 : STD_LOGIC;
    SIGNAL S1478 : STD_LOGIC;
    SIGNAL S1479 : STD_LOGIC;
    SIGNAL S1480 : STD_LOGIC;
    SIGNAL S1481 : STD_LOGIC;
    SIGNAL S1482 : STD_LOGIC;
    SIGNAL S1483 : STD_LOGIC;
    SIGNAL S1484 : STD_LOGIC;
    SIGNAL S1485 : STD_LOGIC;
    SIGNAL S1486 : STD_LOGIC;
    SIGNAL S1487 : STD_LOGIC;
    SIGNAL S1488 : STD_LOGIC;
    SIGNAL S1489 : STD_LOGIC;
    SIGNAL S1490 : STD_LOGIC;
    SIGNAL S1491 : STD_LOGIC;
    SIGNAL S1492 : STD_LOGIC;
    SIGNAL S1493 : STD_LOGIC;
    SIGNAL S1494 : STD_LOGIC;
    SIGNAL S1495 : STD_LOGIC;
    SIGNAL S1496 : STD_LOGIC;
    SIGNAL S1497 : STD_LOGIC;
    SIGNAL S1498 : STD_LOGIC;
    SIGNAL S1499 : STD_LOGIC;
    SIGNAL S1500 : STD_LOGIC;
    SIGNAL S1501 : STD_LOGIC;
    SIGNAL S1502 : STD_LOGIC;
    SIGNAL S1503 : STD_LOGIC;
    SIGNAL S1504 : STD_LOGIC;
    SIGNAL S1505 : STD_LOGIC;
    SIGNAL S1506 : STD_LOGIC;
    SIGNAL S1507 : STD_LOGIC;
    SIGNAL S1508 : STD_LOGIC;
    SIGNAL S1509 : STD_LOGIC;
    SIGNAL S1510 : STD_LOGIC;
    SIGNAL S1511 : STD_LOGIC;
    SIGNAL S1512 : STD_LOGIC;
    SIGNAL S1513 : STD_LOGIC;
    SIGNAL S1514 : STD_LOGIC;
    SIGNAL S1515 : STD_LOGIC;
    SIGNAL S1516 : STD_LOGIC;
    SIGNAL S1517 : STD_LOGIC;
    SIGNAL S1518 : STD_LOGIC;
    SIGNAL S1519 : STD_LOGIC;
    SIGNAL S1520 : STD_LOGIC;
    SIGNAL S1521 : STD_LOGIC;
    SIGNAL S1522 : STD_LOGIC;
    SIGNAL S1523 : STD_LOGIC;
    SIGNAL S1524 : STD_LOGIC;
    SIGNAL S1525 : STD_LOGIC;
    SIGNAL S1526 : STD_LOGIC;
    SIGNAL S1527 : STD_LOGIC;
    SIGNAL S1528 : STD_LOGIC;
    SIGNAL S1529 : STD_LOGIC;
    SIGNAL S1530 : STD_LOGIC;
    SIGNAL S1531 : STD_LOGIC;
    SIGNAL S1532 : STD_LOGIC;
    SIGNAL S1533 : STD_LOGIC;
    SIGNAL S1534 : STD_LOGIC;
    SIGNAL S1535 : STD_LOGIC;
    SIGNAL S1536 : STD_LOGIC;
    SIGNAL S1537 : STD_LOGIC;
    SIGNAL S1538 : STD_LOGIC;
    SIGNAL S1539 : STD_LOGIC;
    SIGNAL S1540 : STD_LOGIC;
    SIGNAL S1541 : STD_LOGIC;
    SIGNAL S1542 : STD_LOGIC;
    SIGNAL S1543 : STD_LOGIC;
    SIGNAL S1544 : STD_LOGIC;
    SIGNAL S1545 : STD_LOGIC;
    SIGNAL S1546 : STD_LOGIC;
    SIGNAL S1547 : STD_LOGIC;
    SIGNAL S1548 : STD_LOGIC;
    SIGNAL S1549 : STD_LOGIC;
    SIGNAL S1550 : STD_LOGIC;
    SIGNAL S1551 : STD_LOGIC;
    SIGNAL S1552 : STD_LOGIC;
    SIGNAL S1553 : STD_LOGIC;
    SIGNAL S1554 : STD_LOGIC;
    SIGNAL S1555 : STD_LOGIC;
    SIGNAL S1556 : STD_LOGIC;
    SIGNAL S1557 : STD_LOGIC;
    SIGNAL S1558 : STD_LOGIC;
    SIGNAL S1559 : STD_LOGIC;
    SIGNAL S1560 : STD_LOGIC;
    SIGNAL S1561 : STD_LOGIC;
    SIGNAL S1562 : STD_LOGIC;
    SIGNAL S1563 : STD_LOGIC;
    SIGNAL S1564 : STD_LOGIC;
    SIGNAL S1565 : STD_LOGIC;
    SIGNAL S1566 : STD_LOGIC;
    SIGNAL S1567 : STD_LOGIC;
    SIGNAL S1568 : STD_LOGIC;
    SIGNAL S1569 : STD_LOGIC;
    SIGNAL S1570 : STD_LOGIC;
    SIGNAL S1571 : STD_LOGIC;
    SIGNAL S1572 : STD_LOGIC;
    SIGNAL S1573 : STD_LOGIC;
    SIGNAL S1574 : STD_LOGIC;
    SIGNAL S1575 : STD_LOGIC;
    SIGNAL S1576 : STD_LOGIC;
    SIGNAL S1577 : STD_LOGIC;
    SIGNAL S1578 : STD_LOGIC;
    SIGNAL S1579 : STD_LOGIC;
    SIGNAL S1580 : STD_LOGIC;
    SIGNAL S1581 : STD_LOGIC;
    SIGNAL S1582 : STD_LOGIC;
    SIGNAL S1583 : STD_LOGIC;
    SIGNAL S1584 : STD_LOGIC;
    SIGNAL S1585 : STD_LOGIC;
    SIGNAL S1586 : STD_LOGIC;
    SIGNAL S1587 : STD_LOGIC;
    SIGNAL S1588 : STD_LOGIC;
    SIGNAL S1589 : STD_LOGIC;
    SIGNAL S1590 : STD_LOGIC;
    SIGNAL S1591 : STD_LOGIC;
    SIGNAL S1592 : STD_LOGIC;
    SIGNAL S1593 : STD_LOGIC;
    SIGNAL S1594 : STD_LOGIC;
    SIGNAL S1595 : STD_LOGIC;
    SIGNAL S1596 : STD_LOGIC;
    SIGNAL S1597 : STD_LOGIC;
    SIGNAL S1598 : STD_LOGIC;
    SIGNAL S1599 : STD_LOGIC;
    SIGNAL S1600 : STD_LOGIC;
    SIGNAL S1601 : STD_LOGIC;
    SIGNAL S1602 : STD_LOGIC;
    SIGNAL S1603 : STD_LOGIC;
    SIGNAL S1604 : STD_LOGIC;
    SIGNAL S1605 : STD_LOGIC;
    SIGNAL S1606 : STD_LOGIC;
    SIGNAL S1607 : STD_LOGIC;
    SIGNAL S1608 : STD_LOGIC;
    SIGNAL S1609 : STD_LOGIC;
    SIGNAL S1610 : STD_LOGIC;
    SIGNAL S1611 : STD_LOGIC;
    SIGNAL S1612 : STD_LOGIC;
    SIGNAL S1613 : STD_LOGIC;
    SIGNAL S1614 : STD_LOGIC;
    SIGNAL S1615 : STD_LOGIC;
    SIGNAL S1616 : STD_LOGIC;
    SIGNAL S1617 : STD_LOGIC;
    SIGNAL S1618 : STD_LOGIC;
    SIGNAL S1619 : STD_LOGIC;
    SIGNAL S1620 : STD_LOGIC;
    SIGNAL S1621 : STD_LOGIC;
    SIGNAL S1622 : STD_LOGIC;
    SIGNAL S1623 : STD_LOGIC;
    SIGNAL S1624 : STD_LOGIC;
    SIGNAL S1625 : STD_LOGIC;
    SIGNAL S1626 : STD_LOGIC;
    SIGNAL S1627 : STD_LOGIC;
    SIGNAL S1628 : STD_LOGIC;
    SIGNAL S1629 : STD_LOGIC;
    SIGNAL S1630 : STD_LOGIC;
    SIGNAL S1631 : STD_LOGIC;
    SIGNAL S1632 : STD_LOGIC;
    SIGNAL S1633 : STD_LOGIC;
    SIGNAL S1634 : STD_LOGIC;
    SIGNAL S1635 : STD_LOGIC;
    SIGNAL S1636 : STD_LOGIC;
    SIGNAL S1637 : STD_LOGIC;
    SIGNAL S1638 : STD_LOGIC;
    SIGNAL S1639 : STD_LOGIC;
    SIGNAL S1640 : STD_LOGIC;
    SIGNAL S1641 : STD_LOGIC;
    SIGNAL S1642 : STD_LOGIC;
    SIGNAL S1643 : STD_LOGIC;
    SIGNAL S1644 : STD_LOGIC;
    SIGNAL S1645 : STD_LOGIC;
    SIGNAL S1646 : STD_LOGIC;
    SIGNAL S1647 : STD_LOGIC;
    SIGNAL S1648 : STD_LOGIC;
    SIGNAL S1649 : STD_LOGIC;
    SIGNAL S1650 : STD_LOGIC;
    SIGNAL S1651 : STD_LOGIC;
    SIGNAL S1652 : STD_LOGIC;
    SIGNAL S1653 : STD_LOGIC;
    SIGNAL S1654 : STD_LOGIC;
    SIGNAL S1655 : STD_LOGIC;
    SIGNAL S1656 : STD_LOGIC;
    SIGNAL S1657 : STD_LOGIC;
    SIGNAL S1658 : STD_LOGIC;
    SIGNAL S1659 : STD_LOGIC;
    SIGNAL S1660 : STD_LOGIC;
    SIGNAL S1661 : STD_LOGIC;
    SIGNAL S1662 : STD_LOGIC;
    SIGNAL S1663 : STD_LOGIC;
    SIGNAL S1664 : STD_LOGIC;
    SIGNAL S1665 : STD_LOGIC;
    SIGNAL S1666 : STD_LOGIC;
    SIGNAL S1667 : STD_LOGIC;
    SIGNAL S1668 : STD_LOGIC;
    SIGNAL S1669 : STD_LOGIC;
    SIGNAL S1670 : STD_LOGIC;
    SIGNAL S1671 : STD_LOGIC;
    SIGNAL S1672 : STD_LOGIC;
    SIGNAL S1673 : STD_LOGIC;
    SIGNAL S1674 : STD_LOGIC;
    SIGNAL S1675 : STD_LOGIC;
    SIGNAL S1676 : STD_LOGIC;
    SIGNAL S1677 : STD_LOGIC;
    SIGNAL S1678 : STD_LOGIC;
    SIGNAL S1679 : STD_LOGIC;
    SIGNAL S1680 : STD_LOGIC;
    SIGNAL S1681 : STD_LOGIC;
    SIGNAL S1682 : STD_LOGIC;
    SIGNAL S1683 : STD_LOGIC;
    SIGNAL S1684 : STD_LOGIC;
    SIGNAL S1685 : STD_LOGIC;
    SIGNAL S1686 : STD_LOGIC;
    SIGNAL S1687 : STD_LOGIC;
    SIGNAL S1688 : STD_LOGIC;
    SIGNAL S1689 : STD_LOGIC;
    SIGNAL S1690 : STD_LOGIC;
    SIGNAL S1691 : STD_LOGIC;
    SIGNAL S1692 : STD_LOGIC;
    SIGNAL S1693 : STD_LOGIC;
    SIGNAL S1694 : STD_LOGIC;
    SIGNAL S1695 : STD_LOGIC;
    SIGNAL S1696 : STD_LOGIC;
    SIGNAL S1697 : STD_LOGIC;
    SIGNAL S1698 : STD_LOGIC;
    SIGNAL S1699 : STD_LOGIC;
    SIGNAL S1700 : STD_LOGIC;
    SIGNAL S1701 : STD_LOGIC;
    SIGNAL S1702 : STD_LOGIC;
    SIGNAL S1703 : STD_LOGIC;
    SIGNAL S1704 : STD_LOGIC;
    SIGNAL S1705 : STD_LOGIC;
    SIGNAL S1706 : STD_LOGIC;
    SIGNAL S1707 : STD_LOGIC;
    SIGNAL S1708 : STD_LOGIC;
    SIGNAL S1709 : STD_LOGIC;
    SIGNAL S1710 : STD_LOGIC;
    SIGNAL S1711 : STD_LOGIC;
    SIGNAL S1712 : STD_LOGIC;
    SIGNAL S1713 : STD_LOGIC;
    SIGNAL S1714 : STD_LOGIC;
    SIGNAL S1715 : STD_LOGIC;
    SIGNAL S1716 : STD_LOGIC;
    SIGNAL S1717 : STD_LOGIC;
    SIGNAL S1718 : STD_LOGIC;
    SIGNAL S1719 : STD_LOGIC;
    SIGNAL S1720 : STD_LOGIC;
    SIGNAL S1721 : STD_LOGIC;
    SIGNAL S1722 : STD_LOGIC;
    SIGNAL S1723 : STD_LOGIC;
    SIGNAL S1724 : STD_LOGIC;
    SIGNAL S1725 : STD_LOGIC;
    SIGNAL S1726 : STD_LOGIC;
    SIGNAL S1727 : STD_LOGIC;
    SIGNAL S1728 : STD_LOGIC;
    SIGNAL S1729 : STD_LOGIC;
    SIGNAL S1730 : STD_LOGIC;
    SIGNAL S1731 : STD_LOGIC;
    SIGNAL S1732 : STD_LOGIC;
    SIGNAL S1733 : STD_LOGIC;
    SIGNAL S1734 : STD_LOGIC;
    SIGNAL S1735 : STD_LOGIC;
    SIGNAL S1736 : STD_LOGIC;
    SIGNAL S1737 : STD_LOGIC;
    SIGNAL S1738 : STD_LOGIC;
    SIGNAL S1739 : STD_LOGIC;
    SIGNAL S1740 : STD_LOGIC;
    SIGNAL S1741 : STD_LOGIC;
    SIGNAL S1742 : STD_LOGIC;
    SIGNAL S1743 : STD_LOGIC;
    SIGNAL S1744 : STD_LOGIC;
    SIGNAL S1745 : STD_LOGIC;
    SIGNAL S1746 : STD_LOGIC;
    SIGNAL S1747 : STD_LOGIC;
    SIGNAL S1748 : STD_LOGIC;
    SIGNAL S1749 : STD_LOGIC;
    SIGNAL S1750 : STD_LOGIC;
    SIGNAL S1751 : STD_LOGIC;
    SIGNAL S1752 : STD_LOGIC;
    SIGNAL S1753 : STD_LOGIC;
    SIGNAL S1754 : STD_LOGIC;
    SIGNAL S1755 : STD_LOGIC;
    SIGNAL S1756 : STD_LOGIC;
    SIGNAL S1757 : STD_LOGIC;
    SIGNAL S1758 : STD_LOGIC;
    SIGNAL S1759 : STD_LOGIC;
    SIGNAL S1760 : STD_LOGIC;
    SIGNAL S1761 : STD_LOGIC;
    SIGNAL S1762 : STD_LOGIC;
    SIGNAL S1763 : STD_LOGIC;
    SIGNAL S1764 : STD_LOGIC;
    SIGNAL S1765 : STD_LOGIC;
    SIGNAL S1766 : STD_LOGIC;
    SIGNAL S1767 : STD_LOGIC;
    SIGNAL S1768 : STD_LOGIC;
    SIGNAL S1769 : STD_LOGIC;
    SIGNAL S1770 : STD_LOGIC;
    SIGNAL S1771 : STD_LOGIC;
    SIGNAL S1772 : STD_LOGIC;
    SIGNAL S1773 : STD_LOGIC;
    SIGNAL S1774 : STD_LOGIC;
    SIGNAL S1775 : STD_LOGIC;
    SIGNAL S1776 : STD_LOGIC;
    SIGNAL S1777 : STD_LOGIC;
    SIGNAL S1778 : STD_LOGIC;
    SIGNAL S1779 : STD_LOGIC;
    SIGNAL S1780 : STD_LOGIC;
    SIGNAL S1781 : STD_LOGIC;
    SIGNAL S1782 : STD_LOGIC;
    SIGNAL S1783 : STD_LOGIC;
    SIGNAL S1784 : STD_LOGIC;
    SIGNAL S1785 : STD_LOGIC;
    SIGNAL S1786 : STD_LOGIC;
    SIGNAL S1787 : STD_LOGIC;
    SIGNAL S1788 : STD_LOGIC;
    SIGNAL S1789 : STD_LOGIC;
    SIGNAL S1790 : STD_LOGIC;
    SIGNAL S1791 : STD_LOGIC;
    SIGNAL S1792 : STD_LOGIC;
    SIGNAL S1793 : STD_LOGIC;
    SIGNAL S1794 : STD_LOGIC;
    SIGNAL S1795 : STD_LOGIC;
    SIGNAL S1796 : STD_LOGIC;
    SIGNAL S1797 : STD_LOGIC;
    SIGNAL S1798 : STD_LOGIC;
    SIGNAL S1799 : STD_LOGIC;
    SIGNAL S1800 : STD_LOGIC;
    SIGNAL S1801 : STD_LOGIC;
    SIGNAL S1802 : STD_LOGIC;
    SIGNAL S1803 : STD_LOGIC;
    SIGNAL S1804 : STD_LOGIC;
    SIGNAL S1805 : STD_LOGIC;
    SIGNAL S1806 : STD_LOGIC;
    SIGNAL S1807 : STD_LOGIC;
    SIGNAL S1808 : STD_LOGIC;
    SIGNAL S1809 : STD_LOGIC;
    SIGNAL S1810 : STD_LOGIC;
    SIGNAL S1811 : STD_LOGIC;
    SIGNAL S1812 : STD_LOGIC;
    SIGNAL S1813 : STD_LOGIC;
    SIGNAL S1814 : STD_LOGIC;
    SIGNAL S1815 : STD_LOGIC;
    SIGNAL S1816 : STD_LOGIC;
    SIGNAL S1817 : STD_LOGIC;
    SIGNAL S1818 : STD_LOGIC;
    SIGNAL S1819 : STD_LOGIC;
    SIGNAL S1820 : STD_LOGIC;
    SIGNAL S1821 : STD_LOGIC;
    SIGNAL S1822 : STD_LOGIC;
    SIGNAL S1823 : STD_LOGIC;
    SIGNAL S1824 : STD_LOGIC;
    SIGNAL S1825 : STD_LOGIC;
    SIGNAL S1826 : STD_LOGIC;
    SIGNAL S1827 : STD_LOGIC;
    SIGNAL S1828 : STD_LOGIC;
    SIGNAL S1829 : STD_LOGIC;
    SIGNAL S1830 : STD_LOGIC;
    SIGNAL S1831 : STD_LOGIC;
    SIGNAL S1832 : STD_LOGIC;
    SIGNAL S1833 : STD_LOGIC;
    SIGNAL S1834 : STD_LOGIC;
    SIGNAL S1835 : STD_LOGIC;
    SIGNAL S1836 : STD_LOGIC;
    SIGNAL S1837 : STD_LOGIC;
    SIGNAL S1838 : STD_LOGIC;
    SIGNAL S1839 : STD_LOGIC;
    SIGNAL S1840 : STD_LOGIC;
    SIGNAL S1841 : STD_LOGIC;
    SIGNAL S1842 : STD_LOGIC;
    SIGNAL S1843 : STD_LOGIC;
    SIGNAL S1844 : STD_LOGIC;
    SIGNAL S1845 : STD_LOGIC;
    SIGNAL S1846 : STD_LOGIC;
    SIGNAL S1847 : STD_LOGIC;
    SIGNAL S1848 : STD_LOGIC;
    SIGNAL S1849 : STD_LOGIC;
    SIGNAL S1850 : STD_LOGIC;
    SIGNAL S1851 : STD_LOGIC;
    SIGNAL S1852 : STD_LOGIC;
    SIGNAL S1853 : STD_LOGIC;
    SIGNAL S1854 : STD_LOGIC;
    SIGNAL S1855 : STD_LOGIC;
    SIGNAL S1856 : STD_LOGIC;
    SIGNAL S1857 : STD_LOGIC;
    SIGNAL S1858 : STD_LOGIC;
    SIGNAL S1859 : STD_LOGIC;
    SIGNAL S1860 : STD_LOGIC;
    SIGNAL S1861 : STD_LOGIC;
    SIGNAL S1862 : STD_LOGIC;
    SIGNAL S1863 : STD_LOGIC;
    SIGNAL S1864 : STD_LOGIC;
    SIGNAL S1865 : STD_LOGIC;
    SIGNAL S1866 : STD_LOGIC;
    SIGNAL S1867 : STD_LOGIC;
    SIGNAL S1868 : STD_LOGIC;
    SIGNAL S1869 : STD_LOGIC;
    SIGNAL S1870 : STD_LOGIC;
    SIGNAL S1871 : STD_LOGIC;
    SIGNAL S1872 : STD_LOGIC;
    SIGNAL S1873 : STD_LOGIC;
    SIGNAL S1874 : STD_LOGIC;
    SIGNAL S1875 : STD_LOGIC;
    SIGNAL S1876 : STD_LOGIC;
    SIGNAL S1877 : STD_LOGIC;
    SIGNAL S1878 : STD_LOGIC;
    SIGNAL S1879 : STD_LOGIC;
    SIGNAL S1880 : STD_LOGIC;
    SIGNAL S1881 : STD_LOGIC;
    SIGNAL S1882 : STD_LOGIC;
    SIGNAL S1883 : STD_LOGIC;
    SIGNAL S1884 : STD_LOGIC;
    SIGNAL S1885 : STD_LOGIC;
    SIGNAL S1886 : STD_LOGIC;
    SIGNAL S1887 : STD_LOGIC;
    SIGNAL S1888 : STD_LOGIC;
    SIGNAL S1889 : STD_LOGIC;
    SIGNAL S1890 : STD_LOGIC;
    SIGNAL S1891 : STD_LOGIC;
    SIGNAL S1892 : STD_LOGIC;
    SIGNAL S1893 : STD_LOGIC;
    SIGNAL S1894 : STD_LOGIC;
    SIGNAL S1895 : STD_LOGIC;
    SIGNAL S1896 : STD_LOGIC;
    SIGNAL S1897 : STD_LOGIC;
    SIGNAL S1898 : STD_LOGIC;
    SIGNAL S1899 : STD_LOGIC;
    SIGNAL S1900 : STD_LOGIC;
    SIGNAL S1901 : STD_LOGIC;
    SIGNAL S1902 : STD_LOGIC;
    SIGNAL S1903 : STD_LOGIC;
    SIGNAL S1904 : STD_LOGIC;
    SIGNAL S1905 : STD_LOGIC;
    SIGNAL S1906 : STD_LOGIC;
    SIGNAL S1907 : STD_LOGIC;
    SIGNAL S1908 : STD_LOGIC;
    SIGNAL S1909 : STD_LOGIC;
    SIGNAL S1910 : STD_LOGIC;
    SIGNAL S1911 : STD_LOGIC;
    SIGNAL S1912 : STD_LOGIC;
    SIGNAL S1913 : STD_LOGIC;
    SIGNAL S1914 : STD_LOGIC;
    SIGNAL S1915 : STD_LOGIC;
    SIGNAL S1916 : STD_LOGIC;
    SIGNAL S1917 : STD_LOGIC;
    SIGNAL S1918 : STD_LOGIC;
    SIGNAL S1919 : STD_LOGIC;
    SIGNAL S1920 : STD_LOGIC;
    SIGNAL S1921 : STD_LOGIC;
    SIGNAL S1922 : STD_LOGIC;
    SIGNAL S1923 : STD_LOGIC;
    SIGNAL S1924 : STD_LOGIC;
    SIGNAL S1925 : STD_LOGIC;
    SIGNAL S1926 : STD_LOGIC;
    SIGNAL S1927 : STD_LOGIC;
    SIGNAL S1928 : STD_LOGIC;
    SIGNAL S1929 : STD_LOGIC;
    SIGNAL S1930 : STD_LOGIC;
    SIGNAL S1931 : STD_LOGIC;
    SIGNAL S1932 : STD_LOGIC;
    SIGNAL S1933 : STD_LOGIC;
    SIGNAL S1934 : STD_LOGIC;
    SIGNAL S1935 : STD_LOGIC;
    SIGNAL S1936 : STD_LOGIC;
    SIGNAL S1937 : STD_LOGIC;
    SIGNAL S1938 : STD_LOGIC;
    SIGNAL S1939 : STD_LOGIC;
    SIGNAL S1940 : STD_LOGIC;
    SIGNAL S1941 : STD_LOGIC;
    SIGNAL S1942 : STD_LOGIC;
    SIGNAL S1943 : STD_LOGIC;
    SIGNAL S1944 : STD_LOGIC;
    SIGNAL S1945 : STD_LOGIC;
    SIGNAL S1946 : STD_LOGIC;
    SIGNAL S1947 : STD_LOGIC;
    SIGNAL S1948 : STD_LOGIC;
    SIGNAL S1949 : STD_LOGIC;
    SIGNAL S1950 : STD_LOGIC;
    SIGNAL S1951 : STD_LOGIC;
    SIGNAL S1952 : STD_LOGIC;
    SIGNAL S1953 : STD_LOGIC;
    SIGNAL S1954 : STD_LOGIC;
    SIGNAL S1955 : STD_LOGIC;
    SIGNAL S1956 : STD_LOGIC;
    SIGNAL S1957 : STD_LOGIC;
    SIGNAL S1958 : STD_LOGIC;
    SIGNAL S1959 : STD_LOGIC;
    SIGNAL S1960 : STD_LOGIC;
    SIGNAL S1961 : STD_LOGIC;
    SIGNAL S1962 : STD_LOGIC;
    SIGNAL S1963 : STD_LOGIC;
    SIGNAL S1964 : STD_LOGIC;
    SIGNAL S1965 : STD_LOGIC;
    SIGNAL S1966 : STD_LOGIC;
    SIGNAL S1967 : STD_LOGIC;
    SIGNAL S1968 : STD_LOGIC;
    SIGNAL S1969 : STD_LOGIC;
    SIGNAL S1970 : STD_LOGIC;
    SIGNAL S1971 : STD_LOGIC;
    SIGNAL S1972 : STD_LOGIC;
    SIGNAL S1973 : STD_LOGIC;
    SIGNAL S1974 : STD_LOGIC;
    SIGNAL S1975 : STD_LOGIC;
    SIGNAL S1976 : STD_LOGIC;
    SIGNAL S1977 : STD_LOGIC;
    SIGNAL S1978 : STD_LOGIC;
    SIGNAL S1979 : STD_LOGIC;
    SIGNAL S1980 : STD_LOGIC;
    SIGNAL S1981 : STD_LOGIC;
    SIGNAL S1982 : STD_LOGIC;
    SIGNAL S1983 : STD_LOGIC;
    SIGNAL S1984 : STD_LOGIC;
    SIGNAL S1985 : STD_LOGIC;
    SIGNAL S1986 : STD_LOGIC;
    SIGNAL S1987 : STD_LOGIC;
    SIGNAL S1988 : STD_LOGIC;
    SIGNAL S1989 : STD_LOGIC;
    SIGNAL S1990 : STD_LOGIC;
    SIGNAL S1991 : STD_LOGIC;
    SIGNAL S1992 : STD_LOGIC;
    SIGNAL S1993 : STD_LOGIC;
    SIGNAL S1994 : STD_LOGIC;
    SIGNAL S1995 : STD_LOGIC;
    SIGNAL S1996 : STD_LOGIC;
    SIGNAL S1997 : STD_LOGIC;
    SIGNAL S1998 : STD_LOGIC;
    SIGNAL S1999 : STD_LOGIC;
    SIGNAL S2000 : STD_LOGIC;
    SIGNAL S2001 : STD_LOGIC;
    SIGNAL S2002 : STD_LOGIC;
    SIGNAL S2003 : STD_LOGIC;
    SIGNAL S2004 : STD_LOGIC;
    SIGNAL S2005 : STD_LOGIC;
    SIGNAL S2006 : STD_LOGIC;
    SIGNAL S2007 : STD_LOGIC;
    SIGNAL S2008 : STD_LOGIC;
    SIGNAL S2009 : STD_LOGIC;
    SIGNAL S2010 : STD_LOGIC;
    SIGNAL S2011 : STD_LOGIC;
    SIGNAL S2012 : STD_LOGIC;
    SIGNAL S2013 : STD_LOGIC;
    SIGNAL S2014 : STD_LOGIC;
    SIGNAL S2015 : STD_LOGIC;
    SIGNAL S2016 : STD_LOGIC;
    SIGNAL S2017 : STD_LOGIC;
    SIGNAL S2018 : STD_LOGIC;
    SIGNAL S2019 : STD_LOGIC;
    SIGNAL S2020 : STD_LOGIC;
    SIGNAL S2021 : STD_LOGIC;
    SIGNAL S2022 : STD_LOGIC;
    SIGNAL S2023 : STD_LOGIC;
    SIGNAL S2024 : STD_LOGIC;
    SIGNAL S2025 : STD_LOGIC;
    SIGNAL S2026 : STD_LOGIC;
    SIGNAL S2027 : STD_LOGIC;
    SIGNAL S2028 : STD_LOGIC;
    SIGNAL S2029 : STD_LOGIC;
    SIGNAL S2030 : STD_LOGIC;
    SIGNAL S2031 : STD_LOGIC;
    SIGNAL S2032 : STD_LOGIC;
    SIGNAL S2033 : STD_LOGIC;
    SIGNAL S2034 : STD_LOGIC;
    SIGNAL S2035 : STD_LOGIC;
    SIGNAL S2036 : STD_LOGIC;
    SIGNAL S2037 : STD_LOGIC;
    SIGNAL S2038 : STD_LOGIC;
    SIGNAL S2039 : STD_LOGIC;
    SIGNAL S2040 : STD_LOGIC;
    SIGNAL S2041 : STD_LOGIC;
    SIGNAL S2042 : STD_LOGIC;
    SIGNAL S2043 : STD_LOGIC;
    SIGNAL S2044 : STD_LOGIC;
    SIGNAL S2045 : STD_LOGIC;
    SIGNAL S2046 : STD_LOGIC;
    SIGNAL S2047 : STD_LOGIC;
    SIGNAL S2048 : STD_LOGIC;
    SIGNAL S2049 : STD_LOGIC;
    SIGNAL S2050 : STD_LOGIC;
    SIGNAL S2051 : STD_LOGIC;
    SIGNAL S2052 : STD_LOGIC;
    SIGNAL S2053 : STD_LOGIC;
    SIGNAL S2054 : STD_LOGIC;
    SIGNAL S2055 : STD_LOGIC;
    SIGNAL S2056 : STD_LOGIC;
    SIGNAL S2057 : STD_LOGIC;
    SIGNAL S2058 : STD_LOGIC;
    SIGNAL S2059 : STD_LOGIC;
    SIGNAL S2060 : STD_LOGIC;
    SIGNAL S2061 : STD_LOGIC;
    SIGNAL S2062 : STD_LOGIC;
    SIGNAL S2063 : STD_LOGIC;
    SIGNAL S2064 : STD_LOGIC;
    SIGNAL S2065 : STD_LOGIC;
    SIGNAL S2066 : STD_LOGIC;
    SIGNAL S2067 : STD_LOGIC;
    SIGNAL S2068 : STD_LOGIC;
    SIGNAL S2069 : STD_LOGIC;
    SIGNAL S2070 : STD_LOGIC;
    SIGNAL S2071 : STD_LOGIC;
    SIGNAL S2072 : STD_LOGIC;
    SIGNAL S2073 : STD_LOGIC;
    SIGNAL S2074 : STD_LOGIC;
    SIGNAL S2075 : STD_LOGIC;
    SIGNAL S2076 : STD_LOGIC;
    SIGNAL S2077 : STD_LOGIC;
    SIGNAL S2078 : STD_LOGIC;
    SIGNAL S2079 : STD_LOGIC;
    SIGNAL S2080 : STD_LOGIC;
    SIGNAL S2081 : STD_LOGIC;
    SIGNAL S2082 : STD_LOGIC;
    SIGNAL S2083 : STD_LOGIC;
    SIGNAL S2084 : STD_LOGIC;
    SIGNAL S2085 : STD_LOGIC;
    SIGNAL S2086 : STD_LOGIC;
    SIGNAL S2087 : STD_LOGIC;
    SIGNAL S2088 : STD_LOGIC;
    SIGNAL S2089 : STD_LOGIC;
    SIGNAL S2090 : STD_LOGIC;
    SIGNAL S2091 : STD_LOGIC;
    SIGNAL S2092 : STD_LOGIC;
    SIGNAL S2093 : STD_LOGIC;
    SIGNAL S2094 : STD_LOGIC;
    SIGNAL S2095 : STD_LOGIC;
    SIGNAL S2096 : STD_LOGIC;
    SIGNAL S2097 : STD_LOGIC;
    SIGNAL S2098 : STD_LOGIC;
    SIGNAL S2099 : STD_LOGIC;
    SIGNAL S2100 : STD_LOGIC;
    SIGNAL S2101 : STD_LOGIC;
    SIGNAL S2102 : STD_LOGIC;
    SIGNAL S2103 : STD_LOGIC;
    SIGNAL S2104 : STD_LOGIC;
    SIGNAL S2105 : STD_LOGIC;
    SIGNAL S2106 : STD_LOGIC;
    SIGNAL S2107 : STD_LOGIC;
    SIGNAL S2108 : STD_LOGIC;
    SIGNAL S2109 : STD_LOGIC;
    SIGNAL S2110 : STD_LOGIC;
    SIGNAL S2111 : STD_LOGIC;
    SIGNAL S2112 : STD_LOGIC;
    SIGNAL S2113 : STD_LOGIC;
    SIGNAL S2114 : STD_LOGIC;
    SIGNAL S2115 : STD_LOGIC;
    SIGNAL S2116 : STD_LOGIC;
    SIGNAL S2117 : STD_LOGIC;
    SIGNAL S2118 : STD_LOGIC;
    SIGNAL S2119 : STD_LOGIC;
    SIGNAL S2120 : STD_LOGIC;
    SIGNAL S2121 : STD_LOGIC;
    SIGNAL S2122 : STD_LOGIC;
    SIGNAL S2123 : STD_LOGIC;
    SIGNAL S2124 : STD_LOGIC;
    SIGNAL S2125 : STD_LOGIC;
    SIGNAL S2126 : STD_LOGIC;
    SIGNAL S2127 : STD_LOGIC;
    SIGNAL S2128 : STD_LOGIC;
    SIGNAL S2129 : STD_LOGIC;
    SIGNAL S2130 : STD_LOGIC;
    SIGNAL S2131 : STD_LOGIC;
    SIGNAL S2132 : STD_LOGIC;
    SIGNAL S2133 : STD_LOGIC;
    SIGNAL S2134 : STD_LOGIC;
    SIGNAL S2135 : STD_LOGIC;
    SIGNAL S2136 : STD_LOGIC;
    SIGNAL S2137 : STD_LOGIC;
    SIGNAL S2138 : STD_LOGIC;
    SIGNAL S2139 : STD_LOGIC;
    SIGNAL S2140 : STD_LOGIC;
    SIGNAL S2141 : STD_LOGIC;
    SIGNAL S2142 : STD_LOGIC;
    SIGNAL S2143 : STD_LOGIC;
    SIGNAL S2144 : STD_LOGIC;
    SIGNAL S2145 : STD_LOGIC;
    SIGNAL S2146 : STD_LOGIC;
    SIGNAL S2147 : STD_LOGIC;
    SIGNAL S2148 : STD_LOGIC;
    SIGNAL S2149 : STD_LOGIC;
    SIGNAL S2150 : STD_LOGIC;
    SIGNAL S2151 : STD_LOGIC;
    SIGNAL S2152 : STD_LOGIC;
    SIGNAL S2153 : STD_LOGIC;
    SIGNAL S2154 : STD_LOGIC;
    SIGNAL S2155 : STD_LOGIC;
    SIGNAL S2156 : STD_LOGIC;
    SIGNAL S2157 : STD_LOGIC;
    SIGNAL S2158 : STD_LOGIC;
    SIGNAL S2159 : STD_LOGIC;
    SIGNAL S2160 : STD_LOGIC;
    SIGNAL S2161 : STD_LOGIC;
    SIGNAL S2162 : STD_LOGIC;
    SIGNAL S2163 : STD_LOGIC;
    SIGNAL S2164 : STD_LOGIC;
    SIGNAL S2165 : STD_LOGIC;
    SIGNAL S2166 : STD_LOGIC;
    SIGNAL S2167 : STD_LOGIC;
    SIGNAL S2168 : STD_LOGIC;
    SIGNAL S2169 : STD_LOGIC;
    SIGNAL S2170 : STD_LOGIC;
    SIGNAL S2171 : STD_LOGIC;
    SIGNAL S2172 : STD_LOGIC;
    SIGNAL S2173 : STD_LOGIC;
    SIGNAL S2174 : STD_LOGIC;
    SIGNAL S2175 : STD_LOGIC;
    SIGNAL S2176 : STD_LOGIC;
    SIGNAL S2177 : STD_LOGIC;
    SIGNAL S2178 : STD_LOGIC;
    SIGNAL S2179 : STD_LOGIC;
    SIGNAL S2180 : STD_LOGIC;
    SIGNAL S2181 : STD_LOGIC;
    SIGNAL S2182 : STD_LOGIC;
    SIGNAL S2183 : STD_LOGIC;
    SIGNAL S2184 : STD_LOGIC;
    SIGNAL S2185 : STD_LOGIC;
    SIGNAL S2186 : STD_LOGIC;
    SIGNAL S2187 : STD_LOGIC;
    SIGNAL S2188 : STD_LOGIC;
    SIGNAL S2189 : STD_LOGIC;
    SIGNAL S2190 : STD_LOGIC;
    SIGNAL S2191 : STD_LOGIC;
    SIGNAL S2192 : STD_LOGIC;
    SIGNAL S2193 : STD_LOGIC;
    SIGNAL S2194 : STD_LOGIC;
    SIGNAL S2195 : STD_LOGIC;
    SIGNAL S2196 : STD_LOGIC;
    SIGNAL S2197 : STD_LOGIC;
    SIGNAL S2198 : STD_LOGIC;
    SIGNAL S2199 : STD_LOGIC;
    SIGNAL S2200 : STD_LOGIC;
    SIGNAL S2201 : STD_LOGIC;
    SIGNAL S2202 : STD_LOGIC;
    SIGNAL S2203 : STD_LOGIC;
    SIGNAL S2204 : STD_LOGIC;
    SIGNAL S2205 : STD_LOGIC;
    SIGNAL S2206 : STD_LOGIC;
    SIGNAL S2207 : STD_LOGIC;
    SIGNAL S2208 : STD_LOGIC;
    SIGNAL S2209 : STD_LOGIC;
    SIGNAL S2210 : STD_LOGIC;
    SIGNAL S2211 : STD_LOGIC;
    SIGNAL S2212 : STD_LOGIC;
    SIGNAL S2213 : STD_LOGIC;
    SIGNAL S2214 : STD_LOGIC;
    SIGNAL S2215 : STD_LOGIC;
    SIGNAL S2216 : STD_LOGIC;
    SIGNAL S2217 : STD_LOGIC;
    SIGNAL S2218 : STD_LOGIC;
    SIGNAL S2219 : STD_LOGIC;
    SIGNAL S2220 : STD_LOGIC;
    SIGNAL S2221 : STD_LOGIC;
    SIGNAL S2222 : STD_LOGIC;
    SIGNAL S2223 : STD_LOGIC;
    SIGNAL S2224 : STD_LOGIC;
    SIGNAL S2225 : STD_LOGIC;
    SIGNAL S2226 : STD_LOGIC;
    SIGNAL S2227 : STD_LOGIC;
    SIGNAL S2228 : STD_LOGIC;
    SIGNAL S2229 : STD_LOGIC;
    SIGNAL S2230 : STD_LOGIC;
    SIGNAL S2231 : STD_LOGIC;
    SIGNAL S2232 : STD_LOGIC;
    SIGNAL S2233 : STD_LOGIC;
    SIGNAL S2234 : STD_LOGIC;
    SIGNAL S2235 : STD_LOGIC;
    SIGNAL S2236 : STD_LOGIC;
    SIGNAL S2237 : STD_LOGIC;
    SIGNAL S2238 : STD_LOGIC;
    SIGNAL S2239 : STD_LOGIC;
    SIGNAL S2240 : STD_LOGIC;
    SIGNAL S2241 : STD_LOGIC;
    SIGNAL S2242 : STD_LOGIC;
    SIGNAL S2243 : STD_LOGIC;
    SIGNAL S2244 : STD_LOGIC;
    SIGNAL S2245 : STD_LOGIC;
    SIGNAL S2246 : STD_LOGIC;
    SIGNAL S2247 : STD_LOGIC;
    SIGNAL S2248 : STD_LOGIC;
    SIGNAL S2249 : STD_LOGIC;
    SIGNAL S2250 : STD_LOGIC;
    SIGNAL S2251 : STD_LOGIC;
    SIGNAL S2252 : STD_LOGIC;
    SIGNAL S2253 : STD_LOGIC;
    SIGNAL S2254 : STD_LOGIC;
    SIGNAL S2255 : STD_LOGIC;
    SIGNAL S2256 : STD_LOGIC;
    SIGNAL S2257 : STD_LOGIC;
    SIGNAL S2258 : STD_LOGIC;
    SIGNAL S2259 : STD_LOGIC;
    SIGNAL S2260 : STD_LOGIC;
    SIGNAL S2261 : STD_LOGIC;
    SIGNAL S2262 : STD_LOGIC;
    SIGNAL S2263 : STD_LOGIC;
    SIGNAL S2264 : STD_LOGIC;
    SIGNAL S2265 : STD_LOGIC;
    SIGNAL S2266 : STD_LOGIC;
    SIGNAL S2267 : STD_LOGIC;
    SIGNAL S2268 : STD_LOGIC;
    SIGNAL S2269 : STD_LOGIC;
    SIGNAL S2270 : STD_LOGIC;
    SIGNAL S2271 : STD_LOGIC;
    SIGNAL S2272 : STD_LOGIC;
    SIGNAL S2273 : STD_LOGIC;
    SIGNAL S2274 : STD_LOGIC;
    SIGNAL S2275 : STD_LOGIC;
    SIGNAL S2276 : STD_LOGIC;
    SIGNAL S2277 : STD_LOGIC;
    SIGNAL S2278 : STD_LOGIC;
    SIGNAL S2279 : STD_LOGIC;
    SIGNAL S2280 : STD_LOGIC;
    SIGNAL S2281 : STD_LOGIC;
    SIGNAL S2282 : STD_LOGIC;
    SIGNAL S2283 : STD_LOGIC;
    SIGNAL S2284 : STD_LOGIC;
    SIGNAL S2285 : STD_LOGIC;
    SIGNAL S2286 : STD_LOGIC;
    SIGNAL S2287 : STD_LOGIC;
    SIGNAL S2288 : STD_LOGIC;
    SIGNAL S2289 : STD_LOGIC;
    SIGNAL S2290 : STD_LOGIC;
    SIGNAL S2291 : STD_LOGIC;
    SIGNAL S2292 : STD_LOGIC;
    SIGNAL S2293 : STD_LOGIC;
    SIGNAL S2294 : STD_LOGIC;
    SIGNAL S2295 : STD_LOGIC;
    SIGNAL S2296 : STD_LOGIC;
    SIGNAL S2297 : STD_LOGIC;
    SIGNAL S2298 : STD_LOGIC;
    SIGNAL S2299 : STD_LOGIC;
    SIGNAL S2300 : STD_LOGIC;
    SIGNAL S2301 : STD_LOGIC;
    SIGNAL S2302 : STD_LOGIC;
    SIGNAL S2303 : STD_LOGIC;
    SIGNAL S2304 : STD_LOGIC;
    SIGNAL S2305 : STD_LOGIC;
    SIGNAL S2306 : STD_LOGIC;
    SIGNAL S2307 : STD_LOGIC;
    SIGNAL S2308 : STD_LOGIC;
    SIGNAL S2309 : STD_LOGIC;
    SIGNAL S2310 : STD_LOGIC;
    SIGNAL S2311 : STD_LOGIC;
    SIGNAL S2312 : STD_LOGIC;
    SIGNAL S2313 : STD_LOGIC;
    SIGNAL S2314 : STD_LOGIC;
    SIGNAL S2315 : STD_LOGIC;
    SIGNAL S2316 : STD_LOGIC;
    SIGNAL S2317 : STD_LOGIC;
    SIGNAL S2318 : STD_LOGIC;
    SIGNAL S2319 : STD_LOGIC;
    SIGNAL S2320 : STD_LOGIC;
    SIGNAL S2321 : STD_LOGIC;
    SIGNAL S2322 : STD_LOGIC;
    SIGNAL S2323 : STD_LOGIC;
    SIGNAL S2324 : STD_LOGIC;
    SIGNAL S2325 : STD_LOGIC;
    SIGNAL S2326 : STD_LOGIC;
    SIGNAL S2327 : STD_LOGIC;
    SIGNAL S2328 : STD_LOGIC;
    SIGNAL S2329 : STD_LOGIC;
    SIGNAL S2330 : STD_LOGIC;
    SIGNAL S2331 : STD_LOGIC;
    SIGNAL S2332 : STD_LOGIC;
    SIGNAL S2333 : STD_LOGIC;
    SIGNAL S2334 : STD_LOGIC;
    SIGNAL S2335 : STD_LOGIC;
    SIGNAL S2336 : STD_LOGIC;
    SIGNAL S2337 : STD_LOGIC;
    SIGNAL S2338 : STD_LOGIC;
    SIGNAL S2339 : STD_LOGIC;
    SIGNAL S2340 : STD_LOGIC;
    SIGNAL S2341 : STD_LOGIC;
    SIGNAL S2342 : STD_LOGIC;
    SIGNAL S2343 : STD_LOGIC;
    SIGNAL S2344 : STD_LOGIC;
    SIGNAL S2345 : STD_LOGIC;
    SIGNAL S2346 : STD_LOGIC;
    SIGNAL S2347 : STD_LOGIC;
    SIGNAL S2348 : STD_LOGIC;
    SIGNAL S2349 : STD_LOGIC;
    SIGNAL S2350 : STD_LOGIC;
    SIGNAL S2351 : STD_LOGIC;
    SIGNAL S2352 : STD_LOGIC;
    SIGNAL S2353 : STD_LOGIC;
    SIGNAL S2354 : STD_LOGIC;
    SIGNAL S2355 : STD_LOGIC;
    SIGNAL S2356 : STD_LOGIC;
    SIGNAL S2357 : STD_LOGIC;
    SIGNAL S2358 : STD_LOGIC;
    SIGNAL S2359 : STD_LOGIC;
    SIGNAL S2360 : STD_LOGIC;
    SIGNAL S2361 : STD_LOGIC;
    SIGNAL S2362 : STD_LOGIC;
    SIGNAL S2363 : STD_LOGIC;
    SIGNAL S2364 : STD_LOGIC;
    SIGNAL S2365 : STD_LOGIC;
    SIGNAL S2366 : STD_LOGIC;
    SIGNAL S2367 : STD_LOGIC;
    SIGNAL S2368 : STD_LOGIC;
    SIGNAL S2369 : STD_LOGIC;
    SIGNAL S2370 : STD_LOGIC;
    SIGNAL S2371 : STD_LOGIC;
    SIGNAL S2372 : STD_LOGIC;
    SIGNAL S2373 : STD_LOGIC;
    SIGNAL S2374 : STD_LOGIC;
    SIGNAL S2375 : STD_LOGIC;
    SIGNAL S2376 : STD_LOGIC;
    SIGNAL S2377 : STD_LOGIC;
    SIGNAL S2378 : STD_LOGIC;
    SIGNAL S2379 : STD_LOGIC;
    SIGNAL S2380 : STD_LOGIC;
    SIGNAL S2381 : STD_LOGIC;
    SIGNAL S2382 : STD_LOGIC;
    SIGNAL S2383 : STD_LOGIC;
    SIGNAL S2384 : STD_LOGIC;
    SIGNAL S2385 : STD_LOGIC;
    SIGNAL S2386 : STD_LOGIC;
    SIGNAL S2387 : STD_LOGIC;
    SIGNAL S2388 : STD_LOGIC;
    SIGNAL S2389 : STD_LOGIC;
    SIGNAL S2390 : STD_LOGIC;
    SIGNAL S2391 : STD_LOGIC;
    SIGNAL S2392 : STD_LOGIC;
    SIGNAL S2393 : STD_LOGIC;
    SIGNAL S2394 : STD_LOGIC;
    SIGNAL S2395 : STD_LOGIC;
    SIGNAL S2396 : STD_LOGIC;
    SIGNAL S2397 : STD_LOGIC;
    SIGNAL S2398 : STD_LOGIC;
    SIGNAL S2399 : STD_LOGIC;
    SIGNAL S2400 : STD_LOGIC;
    SIGNAL S2401 : STD_LOGIC;
    SIGNAL S2402 : STD_LOGIC;
    SIGNAL S2403 : STD_LOGIC;
    SIGNAL S2404 : STD_LOGIC;
    SIGNAL S2405 : STD_LOGIC;
    SIGNAL S2406 : STD_LOGIC;
    SIGNAL S2407 : STD_LOGIC;
    SIGNAL S2408 : STD_LOGIC;
    SIGNAL S2409 : STD_LOGIC;
    SIGNAL S2410 : STD_LOGIC;
    SIGNAL S2411 : STD_LOGIC;
    SIGNAL S2412 : STD_LOGIC;
    SIGNAL S2413 : STD_LOGIC;
    SIGNAL S2414 : STD_LOGIC;
    SIGNAL S2415 : STD_LOGIC;
    SIGNAL S2416 : STD_LOGIC;
    SIGNAL S2417 : STD_LOGIC;
    SIGNAL S2418 : STD_LOGIC;
    SIGNAL S2419 : STD_LOGIC;
    SIGNAL S2420 : STD_LOGIC;
    SIGNAL S2421 : STD_LOGIC;
    SIGNAL S2422 : STD_LOGIC;
    SIGNAL S2423 : STD_LOGIC;
    SIGNAL S2424 : STD_LOGIC;
    SIGNAL S2425 : STD_LOGIC;
    SIGNAL S2426 : STD_LOGIC;
    SIGNAL S2427 : STD_LOGIC;
    SIGNAL S2428 : STD_LOGIC;
    SIGNAL S2429 : STD_LOGIC;
    SIGNAL S2430 : STD_LOGIC;
    SIGNAL S2431 : STD_LOGIC;
    SIGNAL S2432 : STD_LOGIC;
    SIGNAL S2433 : STD_LOGIC;
    SIGNAL S2434 : STD_LOGIC;
    SIGNAL S2435 : STD_LOGIC;
    SIGNAL S2436 : STD_LOGIC;
    SIGNAL S2437 : STD_LOGIC;
    SIGNAL S2438 : STD_LOGIC;
    SIGNAL S2439 : STD_LOGIC;
    SIGNAL S2440 : STD_LOGIC;
    SIGNAL S2441 : STD_LOGIC;
    SIGNAL S2442 : STD_LOGIC;
    SIGNAL S2443 : STD_LOGIC;
    SIGNAL S2444 : STD_LOGIC;
    SIGNAL S2445 : STD_LOGIC;
    SIGNAL S2446 : STD_LOGIC;
    SIGNAL S2447 : STD_LOGIC;
    SIGNAL S2448 : STD_LOGIC;
    SIGNAL S2449 : STD_LOGIC;
    SIGNAL S2450 : STD_LOGIC;
    SIGNAL S2451 : STD_LOGIC;
    SIGNAL S2452 : STD_LOGIC;
    SIGNAL S2453 : STD_LOGIC;
    SIGNAL S2454 : STD_LOGIC;
    SIGNAL S2455 : STD_LOGIC;
    SIGNAL S2456 : STD_LOGIC;
    SIGNAL S2457 : STD_LOGIC;
    SIGNAL S2458 : STD_LOGIC;
    SIGNAL S2459 : STD_LOGIC;
    SIGNAL S2460 : STD_LOGIC;
    SIGNAL S2461 : STD_LOGIC;
    SIGNAL S2462 : STD_LOGIC;
    SIGNAL S2463 : STD_LOGIC;
    SIGNAL S2464 : STD_LOGIC;
    SIGNAL S2465 : STD_LOGIC;
    SIGNAL S2466 : STD_LOGIC;
    SIGNAL S2467 : STD_LOGIC;
    SIGNAL S2468 : STD_LOGIC;
    SIGNAL S2469 : STD_LOGIC;
    SIGNAL S2470 : STD_LOGIC;
    SIGNAL S2471 : STD_LOGIC;
    SIGNAL S2472 : STD_LOGIC;
    SIGNAL S2473 : STD_LOGIC;
    SIGNAL S2474 : STD_LOGIC;
    SIGNAL S2475 : STD_LOGIC;
    SIGNAL S2476 : STD_LOGIC;
    SIGNAL S2477 : STD_LOGIC;
    SIGNAL S2478 : STD_LOGIC;
    SIGNAL S2479 : STD_LOGIC;
    SIGNAL S2480 : STD_LOGIC;
    SIGNAL S2481 : STD_LOGIC;
    SIGNAL S2482 : STD_LOGIC;
    SIGNAL S2483 : STD_LOGIC;
    SIGNAL S2484 : STD_LOGIC;
    SIGNAL S2485 : STD_LOGIC;
    SIGNAL S2486 : STD_LOGIC;
    SIGNAL S2487 : STD_LOGIC;
    SIGNAL S2488 : STD_LOGIC;
    SIGNAL S2489 : STD_LOGIC;
    SIGNAL S2490 : STD_LOGIC;
    SIGNAL S2491 : STD_LOGIC;
    SIGNAL S2492 : STD_LOGIC;
    SIGNAL S2493 : STD_LOGIC;
    SIGNAL S2494 : STD_LOGIC;
    SIGNAL S2495 : STD_LOGIC;
    SIGNAL S2496 : STD_LOGIC;
    SIGNAL S2497 : STD_LOGIC;
    SIGNAL S2498 : STD_LOGIC;
    SIGNAL S2499 : STD_LOGIC;
    SIGNAL S2500 : STD_LOGIC;
    SIGNAL S2501 : STD_LOGIC;
    SIGNAL S2502 : STD_LOGIC;
    SIGNAL S2503 : STD_LOGIC;
    SIGNAL S2504 : STD_LOGIC;
    SIGNAL S2505 : STD_LOGIC;
    SIGNAL S2506 : STD_LOGIC;
    SIGNAL S2507 : STD_LOGIC;
    SIGNAL S2508 : STD_LOGIC;
    SIGNAL S2509 : STD_LOGIC;
    SIGNAL S2510 : STD_LOGIC;
    SIGNAL S2511 : STD_LOGIC;
    SIGNAL S2512 : STD_LOGIC;
    SIGNAL S2513 : STD_LOGIC;
    SIGNAL S2514 : STD_LOGIC;
    SIGNAL S2515 : STD_LOGIC;
    SIGNAL S2516 : STD_LOGIC;
    SIGNAL S2517 : STD_LOGIC;
    SIGNAL S2518 : STD_LOGIC;
    SIGNAL S2519 : STD_LOGIC;
    SIGNAL S2520 : STD_LOGIC;
    SIGNAL S2521 : STD_LOGIC;
    SIGNAL S2522 : STD_LOGIC;
    SIGNAL S2523 : STD_LOGIC;
    SIGNAL S2524 : STD_LOGIC;
    SIGNAL S2525 : STD_LOGIC;
    SIGNAL S2526 : STD_LOGIC;
    SIGNAL S2527 : STD_LOGIC;
    SIGNAL S2528 : STD_LOGIC;
    SIGNAL S2529 : STD_LOGIC;
    SIGNAL S2530 : STD_LOGIC;
    SIGNAL S2531 : STD_LOGIC;
    SIGNAL S2532 : STD_LOGIC;
    SIGNAL S2533 : STD_LOGIC;
    SIGNAL S2534 : STD_LOGIC;
    SIGNAL S2535 : STD_LOGIC;
    SIGNAL S2536 : STD_LOGIC;
    SIGNAL S2537 : STD_LOGIC;
    SIGNAL S2538 : STD_LOGIC;
    SIGNAL S2539 : STD_LOGIC;
    SIGNAL S2540 : STD_LOGIC;
    SIGNAL S2541 : STD_LOGIC;
    SIGNAL S2542 : STD_LOGIC;
    SIGNAL S2543 : STD_LOGIC;
    SIGNAL S2544 : STD_LOGIC;
    SIGNAL S2545 : STD_LOGIC;
    SIGNAL S2546 : STD_LOGIC;
    SIGNAL S2547 : STD_LOGIC;
    SIGNAL S2548 : STD_LOGIC;
    SIGNAL S2549 : STD_LOGIC;
    SIGNAL S2550 : STD_LOGIC;
    SIGNAL S2551 : STD_LOGIC;
    SIGNAL S2552 : STD_LOGIC;
    SIGNAL S2553 : STD_LOGIC;
    SIGNAL S2554 : STD_LOGIC;
    SIGNAL S2555 : STD_LOGIC;
    SIGNAL S2556 : STD_LOGIC;
    SIGNAL S2557 : STD_LOGIC;
    SIGNAL S2558 : STD_LOGIC;
    SIGNAL S2559 : STD_LOGIC;
    SIGNAL S2560 : STD_LOGIC;
    SIGNAL S2561 : STD_LOGIC;
    SIGNAL S2562 : STD_LOGIC;
    SIGNAL S2563 : STD_LOGIC;
    SIGNAL S2564 : STD_LOGIC;
    SIGNAL S2565 : STD_LOGIC;
    SIGNAL S2566 : STD_LOGIC;
    SIGNAL S2567 : STD_LOGIC;
    SIGNAL S2568 : STD_LOGIC;
    SIGNAL S2569 : STD_LOGIC;
    SIGNAL S2570 : STD_LOGIC;
    SIGNAL S2571 : STD_LOGIC;
    SIGNAL S2572 : STD_LOGIC;
    SIGNAL S2573 : STD_LOGIC;
    SIGNAL S2574 : STD_LOGIC;
    SIGNAL S2575 : STD_LOGIC;
    SIGNAL S2576 : STD_LOGIC;
    SIGNAL S2577 : STD_LOGIC;
    SIGNAL S2578 : STD_LOGIC;
    SIGNAL S2579 : STD_LOGIC;
    SIGNAL S2580 : STD_LOGIC;
    SIGNAL S2581 : STD_LOGIC;
    SIGNAL S2582 : STD_LOGIC;
    SIGNAL S2583 : STD_LOGIC;
    SIGNAL S2584 : STD_LOGIC;
    SIGNAL S2585 : STD_LOGIC;
    SIGNAL S2586 : STD_LOGIC;
    SIGNAL S2587 : STD_LOGIC;
    SIGNAL S2588 : STD_LOGIC;
    SIGNAL S2589 : STD_LOGIC;
    SIGNAL S2590 : STD_LOGIC;
    SIGNAL S2591 : STD_LOGIC;
    SIGNAL S2592 : STD_LOGIC;
    SIGNAL S2593 : STD_LOGIC;
    SIGNAL S2594 : STD_LOGIC;
    SIGNAL S2595 : STD_LOGIC;
    SIGNAL S2596 : STD_LOGIC;
    SIGNAL S2597 : STD_LOGIC;
    SIGNAL S2598 : STD_LOGIC;
    SIGNAL S2599 : STD_LOGIC;
    SIGNAL S2600 : STD_LOGIC;
    SIGNAL S2601 : STD_LOGIC;
    SIGNAL S2602 : STD_LOGIC;
    SIGNAL S2603 : STD_LOGIC;
    SIGNAL S2604 : STD_LOGIC;
    SIGNAL S2605 : STD_LOGIC;
    SIGNAL S2606 : STD_LOGIC;
    SIGNAL S2607 : STD_LOGIC;
    SIGNAL S2608 : STD_LOGIC;
    SIGNAL S2609 : STD_LOGIC;
    SIGNAL S2610 : STD_LOGIC;
    SIGNAL S2611 : STD_LOGIC;
    SIGNAL S2612 : STD_LOGIC;
    SIGNAL S2613 : STD_LOGIC;
    SIGNAL S2614 : STD_LOGIC;
    SIGNAL S2615 : STD_LOGIC;
    SIGNAL S2616 : STD_LOGIC;
    SIGNAL S2617 : STD_LOGIC;
    SIGNAL S2618 : STD_LOGIC;
    SIGNAL S2619 : STD_LOGIC;
    SIGNAL S2620 : STD_LOGIC;
    SIGNAL S2621 : STD_LOGIC;
    SIGNAL S2622 : STD_LOGIC;
    SIGNAL S2623 : STD_LOGIC;
    SIGNAL S2624 : STD_LOGIC;
    SIGNAL S2625 : STD_LOGIC;
    SIGNAL S2626 : STD_LOGIC;
    SIGNAL S2627 : STD_LOGIC;
    SIGNAL S2628 : STD_LOGIC;
    SIGNAL S2629 : STD_LOGIC;
    SIGNAL S2630 : STD_LOGIC;
    SIGNAL S2631 : STD_LOGIC;
    SIGNAL S2632 : STD_LOGIC;
    SIGNAL S2633 : STD_LOGIC;
    SIGNAL S2634 : STD_LOGIC;
    SIGNAL S2635 : STD_LOGIC;
    SIGNAL S2636 : STD_LOGIC;
    SIGNAL S2637 : STD_LOGIC;
    SIGNAL S2638 : STD_LOGIC;
    SIGNAL S2639 : STD_LOGIC;
    SIGNAL S2640 : STD_LOGIC;
    SIGNAL S2641 : STD_LOGIC;
    SIGNAL S2642 : STD_LOGIC;
    SIGNAL S2643 : STD_LOGIC;
    SIGNAL S2644 : STD_LOGIC;
    SIGNAL S2645 : STD_LOGIC;
    SIGNAL S2646 : STD_LOGIC;
    SIGNAL S2647 : STD_LOGIC;
    SIGNAL S2648 : STD_LOGIC;
    SIGNAL S2649 : STD_LOGIC;
    SIGNAL S2650 : STD_LOGIC;
    SIGNAL S2651 : STD_LOGIC;
    SIGNAL S2652 : STD_LOGIC;
    SIGNAL S2653 : STD_LOGIC;
    SIGNAL S2654 : STD_LOGIC;
    SIGNAL S2655 : STD_LOGIC;
    SIGNAL S2656 : STD_LOGIC;
    SIGNAL S2657 : STD_LOGIC;
    SIGNAL S2658 : STD_LOGIC;
    SIGNAL S2659 : STD_LOGIC;
    SIGNAL S2660 : STD_LOGIC;
    SIGNAL S2661 : STD_LOGIC;
    SIGNAL S2662 : STD_LOGIC;
    SIGNAL S2663 : STD_LOGIC;
    SIGNAL S2664 : STD_LOGIC;
    SIGNAL S2665 : STD_LOGIC;
    SIGNAL S2666 : STD_LOGIC;
    SIGNAL S2667 : STD_LOGIC;
    SIGNAL S2668 : STD_LOGIC;
    SIGNAL S2669 : STD_LOGIC;
    SIGNAL S2670 : STD_LOGIC;
    SIGNAL S2671 : STD_LOGIC;
    SIGNAL S2672 : STD_LOGIC;
    SIGNAL S2673 : STD_LOGIC;
    SIGNAL S2674 : STD_LOGIC;
    SIGNAL S2675 : STD_LOGIC;
    SIGNAL S2676 : STD_LOGIC;
    SIGNAL S2677 : STD_LOGIC;
    SIGNAL S2678 : STD_LOGIC;
    SIGNAL S2679 : STD_LOGIC;
    SIGNAL S2680 : STD_LOGIC;
    SIGNAL S2681 : STD_LOGIC;
    SIGNAL S2682 : STD_LOGIC;
    SIGNAL S2683 : STD_LOGIC;
    SIGNAL S2684 : STD_LOGIC;
    SIGNAL S2685 : STD_LOGIC;
    SIGNAL S2686 : STD_LOGIC;
    SIGNAL S2687 : STD_LOGIC;
    SIGNAL S2688 : STD_LOGIC;
    SIGNAL S2689 : STD_LOGIC;
    SIGNAL S2690 : STD_LOGIC;
    SIGNAL S2691 : STD_LOGIC;
    SIGNAL S2692 : STD_LOGIC;
    SIGNAL S2693 : STD_LOGIC;
    SIGNAL S2694 : STD_LOGIC;
    SIGNAL S2695 : STD_LOGIC;
    SIGNAL S2696 : STD_LOGIC;
    SIGNAL S2697 : STD_LOGIC;
    SIGNAL S2698 : STD_LOGIC;
    SIGNAL S2699 : STD_LOGIC;
    SIGNAL S2700 : STD_LOGIC;
    SIGNAL S2701 : STD_LOGIC;
    SIGNAL S2702 : STD_LOGIC;
    SIGNAL S2703 : STD_LOGIC;
    SIGNAL S2704 : STD_LOGIC;
    SIGNAL S2705 : STD_LOGIC;
    SIGNAL S2706 : STD_LOGIC;
    SIGNAL S2707 : STD_LOGIC;
    SIGNAL S2708 : STD_LOGIC;
    SIGNAL S2709 : STD_LOGIC;
    SIGNAL S2710 : STD_LOGIC;
    SIGNAL S2711 : STD_LOGIC;
    SIGNAL S2712 : STD_LOGIC;
    SIGNAL S2713 : STD_LOGIC;
    SIGNAL S2714 : STD_LOGIC;
    SIGNAL S2715 : STD_LOGIC;
    SIGNAL S2716 : STD_LOGIC;
    SIGNAL S2717 : STD_LOGIC;
    SIGNAL S2718 : STD_LOGIC;
    SIGNAL S2719 : STD_LOGIC;
    SIGNAL S2720 : STD_LOGIC;
    SIGNAL S2721 : STD_LOGIC;
    SIGNAL S2722 : STD_LOGIC;
    SIGNAL S2723 : STD_LOGIC;
    SIGNAL S2724 : STD_LOGIC;
    SIGNAL S2725 : STD_LOGIC;
    SIGNAL S2726 : STD_LOGIC;
    SIGNAL S2727 : STD_LOGIC;
    SIGNAL S2728 : STD_LOGIC;
    SIGNAL S2729 : STD_LOGIC;
    SIGNAL S2730 : STD_LOGIC;
    SIGNAL S2731 : STD_LOGIC;
    SIGNAL S2732 : STD_LOGIC;
    SIGNAL S2733 : STD_LOGIC;
    SIGNAL S2734 : STD_LOGIC;
    SIGNAL S2735 : STD_LOGIC;
    SIGNAL S2736 : STD_LOGIC;
    SIGNAL S2737 : STD_LOGIC;
    SIGNAL S2738 : STD_LOGIC;
    SIGNAL S2739 : STD_LOGIC;
    SIGNAL S2740 : STD_LOGIC;
    SIGNAL S2741 : STD_LOGIC;
    SIGNAL S2742 : STD_LOGIC;
    SIGNAL S2743 : STD_LOGIC;
    SIGNAL S2744 : STD_LOGIC;
    SIGNAL S2745 : STD_LOGIC;
    SIGNAL S2746 : STD_LOGIC;
    SIGNAL S2747 : STD_LOGIC;
    SIGNAL S2748 : STD_LOGIC;
    SIGNAL S2749 : STD_LOGIC;
    SIGNAL S2750 : STD_LOGIC;
    SIGNAL S2751 : STD_LOGIC;
    SIGNAL S2752 : STD_LOGIC;
    SIGNAL S2753 : STD_LOGIC;
    SIGNAL S2754 : STD_LOGIC;
    SIGNAL S2755 : STD_LOGIC;
    SIGNAL S2756 : STD_LOGIC;
    SIGNAL S2757 : STD_LOGIC;
    SIGNAL S2758 : STD_LOGIC;
    SIGNAL S2759 : STD_LOGIC;
    SIGNAL S2760 : STD_LOGIC;
    SIGNAL S2761 : STD_LOGIC;
    SIGNAL S2762 : STD_LOGIC;
    SIGNAL S2763 : STD_LOGIC;
    SIGNAL S2764 : STD_LOGIC;
    SIGNAL S2765 : STD_LOGIC;
    SIGNAL S2766 : STD_LOGIC;
    SIGNAL S2767 : STD_LOGIC;
    SIGNAL S2768 : STD_LOGIC;
    SIGNAL S2769 : STD_LOGIC;
    SIGNAL S2770 : STD_LOGIC;
    SIGNAL S2771 : STD_LOGIC;
    SIGNAL S2772 : STD_LOGIC;
    SIGNAL S2773 : STD_LOGIC;
    SIGNAL S2774 : STD_LOGIC;
    SIGNAL S2775 : STD_LOGIC;
    SIGNAL S2776 : STD_LOGIC;
    SIGNAL S2777 : STD_LOGIC;
    SIGNAL S2778 : STD_LOGIC;
    SIGNAL S2779 : STD_LOGIC;
    SIGNAL S2780 : STD_LOGIC;
    SIGNAL S2781 : STD_LOGIC;
    SIGNAL S2782 : STD_LOGIC;
    SIGNAL S2783 : STD_LOGIC;
    SIGNAL S2784 : STD_LOGIC;
    SIGNAL S2785 : STD_LOGIC;
    SIGNAL S2786 : STD_LOGIC;
    SIGNAL S2787 : STD_LOGIC;
    SIGNAL S2788 : STD_LOGIC;
    SIGNAL S2789 : STD_LOGIC;
    SIGNAL S2790 : STD_LOGIC;
    SIGNAL S2791 : STD_LOGIC;
    SIGNAL S2792 : STD_LOGIC;
    SIGNAL S2793 : STD_LOGIC;
    SIGNAL S2794 : STD_LOGIC;
    SIGNAL S2795 : STD_LOGIC;
    SIGNAL S2796 : STD_LOGIC;
    SIGNAL S2797 : STD_LOGIC;
    SIGNAL S2798 : STD_LOGIC;
    SIGNAL S2799 : STD_LOGIC;
    SIGNAL S2800 : STD_LOGIC;
    SIGNAL S2801 : STD_LOGIC;
    SIGNAL S2802 : STD_LOGIC;
    SIGNAL S2803 : STD_LOGIC;
    SIGNAL S2804 : STD_LOGIC;
    SIGNAL S2805 : STD_LOGIC;
    SIGNAL S2806 : STD_LOGIC;
    SIGNAL S2807 : STD_LOGIC;
    SIGNAL S2808 : STD_LOGIC;
    SIGNAL S2809 : STD_LOGIC;
    SIGNAL S2810 : STD_LOGIC;
    SIGNAL S2811 : STD_LOGIC;
    SIGNAL S2812 : STD_LOGIC;
    SIGNAL S2813 : STD_LOGIC;
    SIGNAL S2814 : STD_LOGIC;
    SIGNAL S2815 : STD_LOGIC;
    SIGNAL S2816 : STD_LOGIC;
    SIGNAL S2817 : STD_LOGIC;
    SIGNAL S2818 : STD_LOGIC;
    SIGNAL S2819 : STD_LOGIC;
    SIGNAL S2820 : STD_LOGIC;
    SIGNAL S2821 : STD_LOGIC;
    SIGNAL S2822 : STD_LOGIC;
    SIGNAL S2823 : STD_LOGIC;
    SIGNAL S2824 : STD_LOGIC;
    SIGNAL S2825 : STD_LOGIC;
    SIGNAL S2826 : STD_LOGIC;
    SIGNAL S2827 : STD_LOGIC;
    SIGNAL S2828 : STD_LOGIC;
    SIGNAL S2829 : STD_LOGIC;
    SIGNAL S2830 : STD_LOGIC;
    SIGNAL S2831 : STD_LOGIC;
    SIGNAL S2832 : STD_LOGIC;
    SIGNAL S2833 : STD_LOGIC;
    SIGNAL S2834 : STD_LOGIC;
    SIGNAL S2835 : STD_LOGIC;
    SIGNAL S2836 : STD_LOGIC;
    SIGNAL S2837 : STD_LOGIC;
    SIGNAL S2838 : STD_LOGIC;
    SIGNAL S2839 : STD_LOGIC;
    SIGNAL S2840 : STD_LOGIC;
    SIGNAL S2841 : STD_LOGIC;
    SIGNAL S2842 : STD_LOGIC;
    SIGNAL S2843 : STD_LOGIC;
    SIGNAL S2844 : STD_LOGIC;
    SIGNAL S2845 : STD_LOGIC;
    SIGNAL S2846 : STD_LOGIC;
    SIGNAL S2847 : STD_LOGIC;
    SIGNAL S2848 : STD_LOGIC;
    SIGNAL S2849 : STD_LOGIC;
    SIGNAL S2850 : STD_LOGIC;
    SIGNAL S2851 : STD_LOGIC;
    SIGNAL S2852 : STD_LOGIC;
    SIGNAL S2853 : STD_LOGIC;
    SIGNAL S2854 : STD_LOGIC;
    SIGNAL S2855 : STD_LOGIC;
    SIGNAL S2856 : STD_LOGIC;
    SIGNAL S2857 : STD_LOGIC;
    SIGNAL S2858 : STD_LOGIC;
    SIGNAL S2859 : STD_LOGIC;
    SIGNAL S2860 : STD_LOGIC;
    SIGNAL S2861 : STD_LOGIC;
    SIGNAL S2862 : STD_LOGIC;
    SIGNAL S2863 : STD_LOGIC;
    SIGNAL S2864 : STD_LOGIC;
    SIGNAL S2865 : STD_LOGIC;
    SIGNAL S2866 : STD_LOGIC;
    SIGNAL S2867 : STD_LOGIC;
    SIGNAL S2868 : STD_LOGIC;
    SIGNAL S2869 : STD_LOGIC;
    SIGNAL S2870 : STD_LOGIC;
    SIGNAL S2871 : STD_LOGIC;
    SIGNAL S2872 : STD_LOGIC;
    SIGNAL S2873 : STD_LOGIC;
    SIGNAL S2874 : STD_LOGIC;
    SIGNAL S2875 : STD_LOGIC;
    SIGNAL S2876 : STD_LOGIC;
    SIGNAL S2877 : STD_LOGIC;
    SIGNAL S2878 : STD_LOGIC;
    SIGNAL S2879 : STD_LOGIC;
    SIGNAL S2880 : STD_LOGIC;
    SIGNAL S2881 : STD_LOGIC;
    SIGNAL S2882 : STD_LOGIC;
    SIGNAL S2883 : STD_LOGIC;
    SIGNAL S2884 : STD_LOGIC;
    SIGNAL S2885 : STD_LOGIC;
    SIGNAL S2886 : STD_LOGIC;
    SIGNAL S2887 : STD_LOGIC;
    SIGNAL S2888 : STD_LOGIC;
    SIGNAL S2889 : STD_LOGIC;
    SIGNAL S2890 : STD_LOGIC;
    SIGNAL S2891 : STD_LOGIC;
    SIGNAL S2892 : STD_LOGIC;
    SIGNAL S2893 : STD_LOGIC;
    SIGNAL S2894 : STD_LOGIC;
    SIGNAL S2895 : STD_LOGIC;
    SIGNAL S2896 : STD_LOGIC;
    SIGNAL S2897 : STD_LOGIC;
    SIGNAL S2898 : STD_LOGIC;
    SIGNAL S2899 : STD_LOGIC;
    SIGNAL S2900 : STD_LOGIC;
    SIGNAL S2901 : STD_LOGIC;
    SIGNAL S2902 : STD_LOGIC;
    SIGNAL S2903 : STD_LOGIC;
    SIGNAL S2904 : STD_LOGIC;
    SIGNAL S2905 : STD_LOGIC;
    SIGNAL S2906 : STD_LOGIC;
    SIGNAL S2907 : STD_LOGIC;
    SIGNAL S2908 : STD_LOGIC;
    SIGNAL S2909 : STD_LOGIC;
    SIGNAL S2910 : STD_LOGIC;
    SIGNAL S2911 : STD_LOGIC;
    SIGNAL S2912 : STD_LOGIC;
    SIGNAL S2913 : STD_LOGIC;
    SIGNAL S2914 : STD_LOGIC;
    SIGNAL S2915 : STD_LOGIC;
    SIGNAL S2916 : STD_LOGIC;
    SIGNAL S2917 : STD_LOGIC;
    SIGNAL S2918 : STD_LOGIC;
    SIGNAL S2919 : STD_LOGIC;
    SIGNAL S2920 : STD_LOGIC;
    SIGNAL S2921 : STD_LOGIC;
    SIGNAL S2922 : STD_LOGIC;
    SIGNAL S2923 : STD_LOGIC;
    SIGNAL S2924 : STD_LOGIC;
    SIGNAL S2925 : STD_LOGIC;
    SIGNAL S2926 : STD_LOGIC;
    SIGNAL S2927 : STD_LOGIC;
    SIGNAL S2928 : STD_LOGIC;
    SIGNAL S2929 : STD_LOGIC;
    SIGNAL S2930 : STD_LOGIC;
    SIGNAL S2931 : STD_LOGIC;
    SIGNAL S2932 : STD_LOGIC;
    SIGNAL S2933 : STD_LOGIC;
    SIGNAL S2934 : STD_LOGIC;
    SIGNAL S2935 : STD_LOGIC;
    SIGNAL S2936 : STD_LOGIC;
    SIGNAL S2937 : STD_LOGIC;
    SIGNAL S2938 : STD_LOGIC;
    SIGNAL S2939 : STD_LOGIC;
    SIGNAL S2940 : STD_LOGIC;
    SIGNAL S2941 : STD_LOGIC;
    SIGNAL S2942 : STD_LOGIC;
    SIGNAL S2943 : STD_LOGIC;
    SIGNAL S2944 : STD_LOGIC;
    SIGNAL S2945 : STD_LOGIC;
    SIGNAL S2946 : STD_LOGIC;
    SIGNAL S2947 : STD_LOGIC;
    SIGNAL S2948 : STD_LOGIC;
    SIGNAL S2949 : STD_LOGIC;
    SIGNAL S2950 : STD_LOGIC;
    SIGNAL S2951 : STD_LOGIC;
    SIGNAL S2952 : STD_LOGIC;
    SIGNAL S2953 : STD_LOGIC;
    SIGNAL S2954 : STD_LOGIC;
    SIGNAL S2955 : STD_LOGIC;
    SIGNAL S2956 : STD_LOGIC;
    SIGNAL S2957 : STD_LOGIC;
    SIGNAL S2958 : STD_LOGIC;
    SIGNAL S2959 : STD_LOGIC;
    SIGNAL S2960 : STD_LOGIC;
    SIGNAL S2961 : STD_LOGIC;
    SIGNAL S2962 : STD_LOGIC;
    SIGNAL S2963 : STD_LOGIC;
    SIGNAL S2964 : STD_LOGIC;
    SIGNAL S2965 : STD_LOGIC;
    SIGNAL S2966 : STD_LOGIC;
    SIGNAL S2967 : STD_LOGIC;
    SIGNAL S2968 : STD_LOGIC;
    SIGNAL S2969 : STD_LOGIC;
    SIGNAL S2970 : STD_LOGIC;
    SIGNAL S2971 : STD_LOGIC;
    SIGNAL S2972 : STD_LOGIC;
    SIGNAL S2973 : STD_LOGIC;
    SIGNAL S2974 : STD_LOGIC;
    SIGNAL S2975 : STD_LOGIC;
    SIGNAL S2976 : STD_LOGIC;
    SIGNAL S2977 : STD_LOGIC;
    SIGNAL S2978 : STD_LOGIC;
    SIGNAL S2979 : STD_LOGIC;
    SIGNAL S2980 : STD_LOGIC;
    SIGNAL S2981 : STD_LOGIC;
    SIGNAL S2982 : STD_LOGIC;
    SIGNAL S2983 : STD_LOGIC;
    SIGNAL S2984 : STD_LOGIC;
    SIGNAL S2985 : STD_LOGIC;
    SIGNAL S2986 : STD_LOGIC;
    SIGNAL S2987 : STD_LOGIC;
    SIGNAL S2988 : STD_LOGIC;
    SIGNAL S2989 : STD_LOGIC;
    SIGNAL S2990 : STD_LOGIC;
    SIGNAL S2991 : STD_LOGIC;
    SIGNAL S2992 : STD_LOGIC;
    SIGNAL S2993 : STD_LOGIC;
    SIGNAL S2994 : STD_LOGIC;
    SIGNAL S2995 : STD_LOGIC;
    SIGNAL S2996 : STD_LOGIC;
    SIGNAL S2997 : STD_LOGIC;
    SIGNAL S2998 : STD_LOGIC;
    SIGNAL S2999 : STD_LOGIC;
    SIGNAL S3000 : STD_LOGIC;
    SIGNAL S3001 : STD_LOGIC;
    SIGNAL S3002 : STD_LOGIC;
    SIGNAL S3003 : STD_LOGIC;
    SIGNAL S3004 : STD_LOGIC;
    SIGNAL S3005 : STD_LOGIC;
    SIGNAL S3006 : STD_LOGIC;
    SIGNAL S3007 : STD_LOGIC;
    SIGNAL S3008 : STD_LOGIC;
    SIGNAL S3009 : STD_LOGIC;
    SIGNAL S3010 : STD_LOGIC;
    SIGNAL S3011 : STD_LOGIC;
    SIGNAL S3012 : STD_LOGIC;
    SIGNAL S3013 : STD_LOGIC;
    SIGNAL S3014 : STD_LOGIC;
    SIGNAL S3015 : STD_LOGIC;
    SIGNAL S3016 : STD_LOGIC;
    SIGNAL S3017 : STD_LOGIC;
    SIGNAL S3018 : STD_LOGIC;
    SIGNAL S3019 : STD_LOGIC;
    SIGNAL S3020 : STD_LOGIC;
    SIGNAL S3021 : STD_LOGIC;
    SIGNAL S3022 : STD_LOGIC;
    SIGNAL S3023 : STD_LOGIC;
    SIGNAL S3024 : STD_LOGIC;
    SIGNAL S3025 : STD_LOGIC;
    SIGNAL S3026 : STD_LOGIC;
    SIGNAL S3027 : STD_LOGIC;
    SIGNAL S3028 : STD_LOGIC;
    SIGNAL S3029 : STD_LOGIC;
    SIGNAL S3030 : STD_LOGIC;
    SIGNAL S3031 : STD_LOGIC;
    SIGNAL S3032 : STD_LOGIC;
    SIGNAL S3033 : STD_LOGIC;
    SIGNAL S3034 : STD_LOGIC;
    SIGNAL S3035 : STD_LOGIC;
    SIGNAL S3036 : STD_LOGIC;
    SIGNAL S3037 : STD_LOGIC;
    SIGNAL S3038 : STD_LOGIC;
    SIGNAL S3039 : STD_LOGIC;
    SIGNAL S3040 : STD_LOGIC;
    SIGNAL S3041 : STD_LOGIC;
    SIGNAL S3042 : STD_LOGIC;
    SIGNAL S3043 : STD_LOGIC;
    SIGNAL S3044 : STD_LOGIC;
    SIGNAL S3045 : STD_LOGIC;
    SIGNAL S3046 : STD_LOGIC;
    SIGNAL S3047 : STD_LOGIC;
    SIGNAL S3048 : STD_LOGIC;
    SIGNAL S3049 : STD_LOGIC;
    SIGNAL S3050 : STD_LOGIC;
    SIGNAL S3051 : STD_LOGIC;
    SIGNAL S3052 : STD_LOGIC;
    SIGNAL S3053 : STD_LOGIC;
    SIGNAL S3054 : STD_LOGIC;
    SIGNAL S3055 : STD_LOGIC;
    SIGNAL S3056 : STD_LOGIC;
    SIGNAL S3057 : STD_LOGIC;
    SIGNAL S3058 : STD_LOGIC;
    SIGNAL S3059 : STD_LOGIC;
    SIGNAL S3060 : STD_LOGIC;
    SIGNAL S3061 : STD_LOGIC;
    SIGNAL S3062 : STD_LOGIC;
    SIGNAL S3063 : STD_LOGIC;
    SIGNAL S3064 : STD_LOGIC;
    SIGNAL S3065 : STD_LOGIC;
    SIGNAL S3066 : STD_LOGIC;
    SIGNAL S3067 : STD_LOGIC;
    SIGNAL S3068 : STD_LOGIC;
    SIGNAL S3069 : STD_LOGIC;
    SIGNAL S3070 : STD_LOGIC;
    SIGNAL S3071 : STD_LOGIC;
    SIGNAL S3072 : STD_LOGIC;
    SIGNAL S3073 : STD_LOGIC;
    SIGNAL S3074 : STD_LOGIC;
    SIGNAL S3075 : STD_LOGIC;
    SIGNAL S3076 : STD_LOGIC;
    SIGNAL S3077 : STD_LOGIC;
    SIGNAL S3078 : STD_LOGIC;
    SIGNAL S3079 : STD_LOGIC;
    SIGNAL S3080 : STD_LOGIC;
    SIGNAL S3081 : STD_LOGIC;
    SIGNAL S3082 : STD_LOGIC;
    SIGNAL S3083 : STD_LOGIC;
    SIGNAL S3084 : STD_LOGIC;
    SIGNAL S3085 : STD_LOGIC;
    SIGNAL S3086 : STD_LOGIC;
    SIGNAL S3087 : STD_LOGIC;
    SIGNAL S3088 : STD_LOGIC;
    SIGNAL S3089 : STD_LOGIC;
    SIGNAL S3090 : STD_LOGIC;
    SIGNAL S3091 : STD_LOGIC;
    SIGNAL S3092 : STD_LOGIC;
    SIGNAL S3093 : STD_LOGIC;
    SIGNAL S3094 : STD_LOGIC;
    SIGNAL S3095 : STD_LOGIC;
    SIGNAL S3096 : STD_LOGIC;
    SIGNAL S3097 : STD_LOGIC;
    SIGNAL S3098 : STD_LOGIC;
    SIGNAL S3099 : STD_LOGIC;
    SIGNAL S3100 : STD_LOGIC;
    SIGNAL S3101 : STD_LOGIC;
    SIGNAL S3102 : STD_LOGIC;
    SIGNAL S3103 : STD_LOGIC;
    SIGNAL S3104 : STD_LOGIC;
    SIGNAL S3105 : STD_LOGIC;
    SIGNAL S3106 : STD_LOGIC;
    SIGNAL S3107 : STD_LOGIC;
    SIGNAL S3108 : STD_LOGIC;
    SIGNAL S3109 : STD_LOGIC;
    SIGNAL S3110 : STD_LOGIC;
    SIGNAL S3111 : STD_LOGIC;
    SIGNAL S3112 : STD_LOGIC;
    SIGNAL S3113 : STD_LOGIC;
    SIGNAL S3114 : STD_LOGIC;
    SIGNAL S3115 : STD_LOGIC;
    SIGNAL S3116 : STD_LOGIC;
    SIGNAL S3117 : STD_LOGIC;
    SIGNAL S3118 : STD_LOGIC;
    SIGNAL S3119 : STD_LOGIC;
    SIGNAL S3120 : STD_LOGIC;
    SIGNAL S3121 : STD_LOGIC;
    SIGNAL S3122 : STD_LOGIC;
    SIGNAL S3123 : STD_LOGIC;
    SIGNAL S3124 : STD_LOGIC;
    SIGNAL S3125 : STD_LOGIC;
    SIGNAL S3126 : STD_LOGIC;
    SIGNAL S3127 : STD_LOGIC;
    SIGNAL S3128 : STD_LOGIC;
    SIGNAL S3129 : STD_LOGIC;
    SIGNAL S3130 : STD_LOGIC;
    SIGNAL S3131 : STD_LOGIC;
    SIGNAL S3132 : STD_LOGIC;
    SIGNAL S3133 : STD_LOGIC;
    SIGNAL S3134 : STD_LOGIC;
    SIGNAL S3135 : STD_LOGIC;
    SIGNAL S3136 : STD_LOGIC;
    SIGNAL S3137 : STD_LOGIC;
    SIGNAL S3138 : STD_LOGIC;
    SIGNAL S3139 : STD_LOGIC;
    SIGNAL S3140 : STD_LOGIC;
    SIGNAL S3141 : STD_LOGIC;
    SIGNAL S3142 : STD_LOGIC;
    SIGNAL S3143 : STD_LOGIC;
    SIGNAL S3144 : STD_LOGIC;
    SIGNAL S3145 : STD_LOGIC;
    SIGNAL S3146 : STD_LOGIC;
    SIGNAL S3147 : STD_LOGIC;
    SIGNAL S3148 : STD_LOGIC;
    SIGNAL S3149 : STD_LOGIC;
    SIGNAL S3150 : STD_LOGIC;
    SIGNAL S3151 : STD_LOGIC;
    SIGNAL S3152 : STD_LOGIC;
    SIGNAL S3153 : STD_LOGIC;
    SIGNAL S3154 : STD_LOGIC;
    SIGNAL S3155 : STD_LOGIC;
    SIGNAL S3156 : STD_LOGIC;
    SIGNAL S3157 : STD_LOGIC;
    SIGNAL S3158 : STD_LOGIC;
    SIGNAL S3159 : STD_LOGIC;
    SIGNAL S3160 : STD_LOGIC;
    SIGNAL S3161 : STD_LOGIC;
    SIGNAL S3162 : STD_LOGIC;
    SIGNAL S3163 : STD_LOGIC;
    SIGNAL S3164 : STD_LOGIC;
    SIGNAL S3165 : STD_LOGIC;
    SIGNAL S3166 : STD_LOGIC;
    SIGNAL S3167 : STD_LOGIC;
    SIGNAL S3168 : STD_LOGIC;
    SIGNAL S3169 : STD_LOGIC;
    SIGNAL S3170 : STD_LOGIC;
    SIGNAL S3171 : STD_LOGIC;
    SIGNAL S3172 : STD_LOGIC;
    SIGNAL S3173 : STD_LOGIC;
    SIGNAL S3174 : STD_LOGIC;
    SIGNAL S3175 : STD_LOGIC;
    SIGNAL S3176 : STD_LOGIC;
    SIGNAL S3177 : STD_LOGIC;
    SIGNAL S3178 : STD_LOGIC;
    SIGNAL S3179 : STD_LOGIC;
    SIGNAL S3180 : STD_LOGIC;
    SIGNAL S3181 : STD_LOGIC;
    SIGNAL S3182 : STD_LOGIC;
    SIGNAL S3183 : STD_LOGIC;
    SIGNAL S3184 : STD_LOGIC;
    SIGNAL S3185 : STD_LOGIC;
    SIGNAL S3186 : STD_LOGIC;
    SIGNAL S3187 : STD_LOGIC;
    SIGNAL S3188 : STD_LOGIC;
    SIGNAL S3189 : STD_LOGIC;
    SIGNAL S3190 : STD_LOGIC;
    SIGNAL S3191 : STD_LOGIC;
    SIGNAL S3192 : STD_LOGIC;
    SIGNAL S3193 : STD_LOGIC;
    SIGNAL S3194 : STD_LOGIC;
    SIGNAL S3195 : STD_LOGIC;
    SIGNAL S3196 : STD_LOGIC;
    SIGNAL S3197 : STD_LOGIC;
    SIGNAL S3198 : STD_LOGIC;
    SIGNAL S3199 : STD_LOGIC;
    SIGNAL S3200 : STD_LOGIC;
    SIGNAL S3201 : STD_LOGIC;
    SIGNAL S3202 : STD_LOGIC;
    SIGNAL S3203 : STD_LOGIC;
    SIGNAL S3204 : STD_LOGIC;
    SIGNAL S3205 : STD_LOGIC;
    SIGNAL S3206 : STD_LOGIC;
    SIGNAL S3207 : STD_LOGIC;
    SIGNAL S3208 : STD_LOGIC;
    SIGNAL S3209 : STD_LOGIC;
    SIGNAL S3210 : STD_LOGIC;
    SIGNAL S3211 : STD_LOGIC;
    SIGNAL S3212 : STD_LOGIC;
    SIGNAL S3213 : STD_LOGIC;
    SIGNAL S3214 : STD_LOGIC;
    SIGNAL S3215 : STD_LOGIC;
    SIGNAL S3216 : STD_LOGIC;
    SIGNAL S3217 : STD_LOGIC;
    SIGNAL S3218 : STD_LOGIC;
    SIGNAL S3219 : STD_LOGIC;
    SIGNAL S3220 : STD_LOGIC;
    SIGNAL S3221 : STD_LOGIC;
    SIGNAL S3222 : STD_LOGIC;
    SIGNAL S3223 : STD_LOGIC;
    SIGNAL S3224 : STD_LOGIC;
    SIGNAL S3225 : STD_LOGIC;
    SIGNAL S3226 : STD_LOGIC;
    SIGNAL S3227 : STD_LOGIC;
    SIGNAL S3228 : STD_LOGIC;
    SIGNAL S3229 : STD_LOGIC;
    SIGNAL S3230 : STD_LOGIC;
    SIGNAL S3231 : STD_LOGIC;
    SIGNAL S3232 : STD_LOGIC;
    SIGNAL S3233 : STD_LOGIC;
    SIGNAL S3234 : STD_LOGIC;
    SIGNAL S3235 : STD_LOGIC;
    SIGNAL S3236 : STD_LOGIC;
    SIGNAL S3237 : STD_LOGIC;
    SIGNAL S3238 : STD_LOGIC;
    SIGNAL S3239 : STD_LOGIC;
    SIGNAL S3240 : STD_LOGIC;
    SIGNAL S3241 : STD_LOGIC;
    SIGNAL S3242 : STD_LOGIC;
    SIGNAL S3243 : STD_LOGIC;
    SIGNAL S3244 : STD_LOGIC;
    SIGNAL S3245 : STD_LOGIC;
    SIGNAL S3246 : STD_LOGIC;
    SIGNAL S3247 : STD_LOGIC;
    SIGNAL S3248 : STD_LOGIC;
    SIGNAL S3249 : STD_LOGIC;
    SIGNAL S3250 : STD_LOGIC;
    SIGNAL S3251 : STD_LOGIC;
    SIGNAL S3252 : STD_LOGIC;
    SIGNAL S3253 : STD_LOGIC;
    SIGNAL S3254 : STD_LOGIC;
    SIGNAL S3255 : STD_LOGIC;
    SIGNAL S3256 : STD_LOGIC;
    SIGNAL S3257 : STD_LOGIC;
    SIGNAL S3258 : STD_LOGIC;
    SIGNAL S3259 : STD_LOGIC;
    SIGNAL S3260 : STD_LOGIC;
    SIGNAL S3261 : STD_LOGIC;
    SIGNAL S3262 : STD_LOGIC;
    SIGNAL S3263 : STD_LOGIC;
    SIGNAL S3264 : STD_LOGIC;
    SIGNAL S3265 : STD_LOGIC;
    SIGNAL S3266 : STD_LOGIC;
    SIGNAL S3267 : STD_LOGIC;
    SIGNAL S3268 : STD_LOGIC;
    SIGNAL S3269 : STD_LOGIC;
    SIGNAL S3270 : STD_LOGIC;
    SIGNAL S3271 : STD_LOGIC;
    SIGNAL S3272 : STD_LOGIC;
    SIGNAL S3273 : STD_LOGIC;
    SIGNAL S3274 : STD_LOGIC;
    SIGNAL S3275 : STD_LOGIC;
    SIGNAL S3276 : STD_LOGIC;
    SIGNAL S3277 : STD_LOGIC;
    SIGNAL S3278 : STD_LOGIC;
    SIGNAL S3279 : STD_LOGIC;
    SIGNAL S3280 : STD_LOGIC;
    SIGNAL S3281 : STD_LOGIC;
    SIGNAL S3282 : STD_LOGIC;
    SIGNAL S3283 : STD_LOGIC;
    SIGNAL S3284 : STD_LOGIC;
    SIGNAL S3285 : STD_LOGIC;
    SIGNAL S3286 : STD_LOGIC;
    SIGNAL S3287 : STD_LOGIC;
    SIGNAL S3288 : STD_LOGIC;
    SIGNAL S3289 : STD_LOGIC;
    SIGNAL S3290 : STD_LOGIC;
    SIGNAL S3291 : STD_LOGIC;
    SIGNAL S3292 : STD_LOGIC;
    SIGNAL S3293 : STD_LOGIC;
    SIGNAL S3294 : STD_LOGIC;
    SIGNAL S3295 : STD_LOGIC;
    SIGNAL S3296 : STD_LOGIC;
    SIGNAL S3297 : STD_LOGIC;
    SIGNAL S3298 : STD_LOGIC;
    SIGNAL S3299 : STD_LOGIC;
    SIGNAL S3300 : STD_LOGIC;
    SIGNAL S3301 : STD_LOGIC;
    SIGNAL S3302 : STD_LOGIC;
    SIGNAL S3303 : STD_LOGIC;
    SIGNAL S3304 : STD_LOGIC;
    SIGNAL S3305 : STD_LOGIC;
    SIGNAL S3306 : STD_LOGIC;
    SIGNAL S3307 : STD_LOGIC;
    SIGNAL S3308 : STD_LOGIC;
    SIGNAL S3309 : STD_LOGIC;
    SIGNAL S3310 : STD_LOGIC;
    SIGNAL S3311 : STD_LOGIC;
    SIGNAL S3312 : STD_LOGIC;
    SIGNAL S3313 : STD_LOGIC;
    SIGNAL S3314 : STD_LOGIC;
    SIGNAL S3315 : STD_LOGIC;
    SIGNAL S3316 : STD_LOGIC;
    SIGNAL S3317 : STD_LOGIC;
    SIGNAL S3318 : STD_LOGIC;
    SIGNAL S3319 : STD_LOGIC;
    SIGNAL S3320 : STD_LOGIC;
    SIGNAL S3321 : STD_LOGIC;
    SIGNAL S3322 : STD_LOGIC;
    SIGNAL S3323 : STD_LOGIC;
    SIGNAL S3324 : STD_LOGIC;
    SIGNAL S3325 : STD_LOGIC;
    SIGNAL S3326 : STD_LOGIC;
    SIGNAL S3327 : STD_LOGIC;
    SIGNAL S3328 : STD_LOGIC;
    SIGNAL S3329 : STD_LOGIC;
    SIGNAL S3330 : STD_LOGIC;
    SIGNAL S3331 : STD_LOGIC;
    SIGNAL S3332 : STD_LOGIC;
    SIGNAL S3333 : STD_LOGIC;
    SIGNAL S3334 : STD_LOGIC;
    SIGNAL S3335 : STD_LOGIC;
    SIGNAL S3336 : STD_LOGIC;
    SIGNAL S3337 : STD_LOGIC;
    SIGNAL S3338 : STD_LOGIC;
    SIGNAL S3339 : STD_LOGIC;
    SIGNAL S3340 : STD_LOGIC;
    SIGNAL S3341 : STD_LOGIC;
    SIGNAL S3342 : STD_LOGIC;
    SIGNAL S3343 : STD_LOGIC;
    SIGNAL S3344 : STD_LOGIC;
    SIGNAL S3345 : STD_LOGIC;
    SIGNAL S3346 : STD_LOGIC;
    SIGNAL S3347 : STD_LOGIC;
    SIGNAL S3348 : STD_LOGIC;
    SIGNAL S3349 : STD_LOGIC;
    SIGNAL S3350 : STD_LOGIC;
    SIGNAL S3351 : STD_LOGIC;
    SIGNAL S3352 : STD_LOGIC;
    SIGNAL S3353 : STD_LOGIC;
    SIGNAL S3354 : STD_LOGIC;
    SIGNAL S3355 : STD_LOGIC;
    SIGNAL S3356 : STD_LOGIC;
    SIGNAL S3357 : STD_LOGIC;
    SIGNAL S3358 : STD_LOGIC;
    SIGNAL S3359 : STD_LOGIC;
    SIGNAL S3360 : STD_LOGIC;
    SIGNAL S3361 : STD_LOGIC;
    SIGNAL S3362 : STD_LOGIC;
    SIGNAL S3363 : STD_LOGIC;
    SIGNAL S3364 : STD_LOGIC;
    SIGNAL S3365 : STD_LOGIC;
    SIGNAL S3366 : STD_LOGIC;
    SIGNAL S3367 : STD_LOGIC;
    SIGNAL S3368 : STD_LOGIC;
    SIGNAL S3369 : STD_LOGIC;
    SIGNAL S3370 : STD_LOGIC;
    SIGNAL S3371 : STD_LOGIC;
    SIGNAL S3372 : STD_LOGIC;
    SIGNAL S3373 : STD_LOGIC;
    SIGNAL S3374 : STD_LOGIC;
    SIGNAL S3375 : STD_LOGIC;
    SIGNAL S3376 : STD_LOGIC;
    SIGNAL S3377 : STD_LOGIC;
    SIGNAL S3378 : STD_LOGIC;
    SIGNAL S3379 : STD_LOGIC;
    SIGNAL S3380 : STD_LOGIC;
    SIGNAL S3381 : STD_LOGIC;
    SIGNAL S3382 : STD_LOGIC;
    SIGNAL S3383 : STD_LOGIC;
    SIGNAL S3384 : STD_LOGIC;
    SIGNAL S3385 : STD_LOGIC;
    SIGNAL S3386 : STD_LOGIC;
    SIGNAL S3387 : STD_LOGIC;
    SIGNAL S3388 : STD_LOGIC;
    SIGNAL S3389 : STD_LOGIC;
    SIGNAL S3390 : STD_LOGIC;
    SIGNAL S3391 : STD_LOGIC;
    SIGNAL S3392 : STD_LOGIC;
    SIGNAL S3393 : STD_LOGIC;
    SIGNAL S3394 : STD_LOGIC;
    SIGNAL S3395 : STD_LOGIC;
    SIGNAL S3396 : STD_LOGIC;
    SIGNAL S3397 : STD_LOGIC;
    SIGNAL S3398 : STD_LOGIC;
    SIGNAL S3399 : STD_LOGIC;
    SIGNAL S3400 : STD_LOGIC;
    SIGNAL S3401 : STD_LOGIC;
    SIGNAL S3402 : STD_LOGIC;
    SIGNAL S3403 : STD_LOGIC;
    SIGNAL S3404 : STD_LOGIC;
    SIGNAL S3405 : STD_LOGIC;
    SIGNAL S3406 : STD_LOGIC;
    SIGNAL S3407 : STD_LOGIC;
    SIGNAL S3408 : STD_LOGIC;
    SIGNAL S3409 : STD_LOGIC;
    SIGNAL S3410 : STD_LOGIC;
    SIGNAL S3411 : STD_LOGIC;
    SIGNAL S3412 : STD_LOGIC;
    SIGNAL S3413 : STD_LOGIC;
    SIGNAL S3414 : STD_LOGIC;
    SIGNAL S3415 : STD_LOGIC;
    SIGNAL S3416 : STD_LOGIC;
    SIGNAL S3417 : STD_LOGIC;
    SIGNAL S3418 : STD_LOGIC;
    SIGNAL S3419 : STD_LOGIC;
    SIGNAL S3420 : STD_LOGIC;
    SIGNAL S3421 : STD_LOGIC;
    SIGNAL S3422 : STD_LOGIC;
    SIGNAL S3423 : STD_LOGIC;
    SIGNAL S3424 : STD_LOGIC;
    SIGNAL S3425 : STD_LOGIC;
    SIGNAL S3426 : STD_LOGIC;
    SIGNAL S3427 : STD_LOGIC;
    SIGNAL S3428 : STD_LOGIC;
    SIGNAL S3429 : STD_LOGIC;
    SIGNAL S3430 : STD_LOGIC;
    SIGNAL S3431 : STD_LOGIC;
    SIGNAL S3432 : STD_LOGIC;
    SIGNAL S3433 : STD_LOGIC;
    SIGNAL S3434 : STD_LOGIC;
    SIGNAL S3435 : STD_LOGIC;
    SIGNAL S3436 : STD_LOGIC;
    SIGNAL S3437 : STD_LOGIC;
    SIGNAL S3438 : STD_LOGIC;
    SIGNAL S3439 : STD_LOGIC;
    SIGNAL S3440 : STD_LOGIC;
    SIGNAL S3441 : STD_LOGIC;
    SIGNAL S3442 : STD_LOGIC;
    SIGNAL S3443 : STD_LOGIC;
    SIGNAL S3444 : STD_LOGIC;
    SIGNAL S3445 : STD_LOGIC;
    SIGNAL S3446 : STD_LOGIC;
    SIGNAL S3447 : STD_LOGIC;
    SIGNAL S3448 : STD_LOGIC;
    SIGNAL S3449 : STD_LOGIC;
    SIGNAL S3450 : STD_LOGIC;
    SIGNAL S3451 : STD_LOGIC;
    SIGNAL S3452 : STD_LOGIC;
    SIGNAL S3453 : STD_LOGIC;
    SIGNAL S3454 : STD_LOGIC;
    SIGNAL S3455 : STD_LOGIC;
    SIGNAL S3456 : STD_LOGIC;
    SIGNAL S3457 : STD_LOGIC;
    SIGNAL S3458 : STD_LOGIC;
    SIGNAL S3459 : STD_LOGIC;
    SIGNAL S3460 : STD_LOGIC;
    SIGNAL S3461 : STD_LOGIC;
    SIGNAL S3462 : STD_LOGIC;
    SIGNAL S3463 : STD_LOGIC;
    SIGNAL S3464 : STD_LOGIC;
    SIGNAL S3465 : STD_LOGIC;
    SIGNAL S3466 : STD_LOGIC;
    SIGNAL S3467 : STD_LOGIC;
    SIGNAL S3468 : STD_LOGIC;
    SIGNAL S3469 : STD_LOGIC;
    SIGNAL S3470 : STD_LOGIC;
    SIGNAL S3471 : STD_LOGIC;
    SIGNAL S3472 : STD_LOGIC;
    SIGNAL S3473 : STD_LOGIC;
    SIGNAL S3474 : STD_LOGIC;
    SIGNAL S3475 : STD_LOGIC;
    SIGNAL S3476 : STD_LOGIC;
    SIGNAL S3477 : STD_LOGIC;
    SIGNAL S3478 : STD_LOGIC;
    SIGNAL S3479 : STD_LOGIC;
    SIGNAL S3480 : STD_LOGIC;
    SIGNAL S3481 : STD_LOGIC;
    SIGNAL S3482 : STD_LOGIC;
    SIGNAL S3483 : STD_LOGIC;
    SIGNAL S3484 : STD_LOGIC;
    SIGNAL S3485 : STD_LOGIC;
    SIGNAL S3486 : STD_LOGIC;
    SIGNAL S3487 : STD_LOGIC;
    SIGNAL S3488 : STD_LOGIC;
    SIGNAL S3489 : STD_LOGIC;
    SIGNAL S3490 : STD_LOGIC;
    SIGNAL S3491 : STD_LOGIC;
    SIGNAL S3492 : STD_LOGIC;
    SIGNAL S3493 : STD_LOGIC;
    SIGNAL S3494 : STD_LOGIC;
    SIGNAL S3495 : STD_LOGIC;
    SIGNAL S3496 : STD_LOGIC;
    SIGNAL S3497 : STD_LOGIC;
    SIGNAL S3498 : STD_LOGIC;
    SIGNAL S3499 : STD_LOGIC;
    SIGNAL S3500 : STD_LOGIC;
    SIGNAL S3501 : STD_LOGIC;
    SIGNAL S3502 : STD_LOGIC;
    SIGNAL S3503 : STD_LOGIC;
    SIGNAL S3504 : STD_LOGIC;
    SIGNAL S3505 : STD_LOGIC;
    SIGNAL S3506 : STD_LOGIC;
    SIGNAL S3507 : STD_LOGIC;
    SIGNAL S3508 : STD_LOGIC;
    SIGNAL S3509 : STD_LOGIC;
    SIGNAL S3510 : STD_LOGIC;
    SIGNAL S3511 : STD_LOGIC;
    SIGNAL S3512 : STD_LOGIC;
    SIGNAL S3513 : STD_LOGIC;
    SIGNAL S3514 : STD_LOGIC;
    SIGNAL S3515 : STD_LOGIC;
    SIGNAL S3516 : STD_LOGIC;
    SIGNAL S3517 : STD_LOGIC;
    SIGNAL S3518 : STD_LOGIC;
    SIGNAL S3519 : STD_LOGIC;
    SIGNAL S3520 : STD_LOGIC;
    SIGNAL S3521 : STD_LOGIC;
    SIGNAL S3522 : STD_LOGIC;
    SIGNAL S3523 : STD_LOGIC;
    SIGNAL S3524 : STD_LOGIC;
    SIGNAL S3525 : STD_LOGIC;
    SIGNAL S3526 : STD_LOGIC;
    SIGNAL S3527 : STD_LOGIC;
    SIGNAL S3528 : STD_LOGIC;
    SIGNAL S3529 : STD_LOGIC;
    SIGNAL S3530 : STD_LOGIC;
    SIGNAL S3531 : STD_LOGIC;
    SIGNAL S3532 : STD_LOGIC;
    SIGNAL S3533 : STD_LOGIC;
    SIGNAL S3534 : STD_LOGIC;
    SIGNAL S3535 : STD_LOGIC;
    SIGNAL S3536 : STD_LOGIC;
    SIGNAL S3537 : STD_LOGIC;
    SIGNAL S3538 : STD_LOGIC;
    SIGNAL S3539 : STD_LOGIC;
    SIGNAL S3540 : STD_LOGIC;
    SIGNAL S3541 : STD_LOGIC;
    SIGNAL S3542 : STD_LOGIC;
    SIGNAL S3543 : STD_LOGIC;
    SIGNAL S3544 : STD_LOGIC;
    SIGNAL S3545 : STD_LOGIC;
    SIGNAL S3546 : STD_LOGIC;
    SIGNAL S3547 : STD_LOGIC;
    SIGNAL S3548 : STD_LOGIC;
    SIGNAL S3549 : STD_LOGIC;
    SIGNAL S3550 : STD_LOGIC;
    SIGNAL S3551 : STD_LOGIC;
    SIGNAL S3552 : STD_LOGIC;
    SIGNAL S3553 : STD_LOGIC;
    SIGNAL S3554 : STD_LOGIC;
    SIGNAL S3555 : STD_LOGIC;
    SIGNAL S3556 : STD_LOGIC;
    SIGNAL S3557 : STD_LOGIC;
    SIGNAL S3558 : STD_LOGIC;
    SIGNAL S3559 : STD_LOGIC;
    SIGNAL S3560 : STD_LOGIC;
    SIGNAL S3561 : STD_LOGIC;
    SIGNAL S3562 : STD_LOGIC;
    SIGNAL S3563 : STD_LOGIC;
    SIGNAL S3564 : STD_LOGIC;
    SIGNAL S3565 : STD_LOGIC;
    SIGNAL S3566 : STD_LOGIC;
    SIGNAL S3567 : STD_LOGIC;
    SIGNAL S3568 : STD_LOGIC;
    SIGNAL S3569 : STD_LOGIC;
    SIGNAL S3570 : STD_LOGIC;
    SIGNAL S3571 : STD_LOGIC;
    SIGNAL S3572 : STD_LOGIC;
    SIGNAL S3573 : STD_LOGIC;
    SIGNAL S3574 : STD_LOGIC;
    SIGNAL S3575 : STD_LOGIC;
    SIGNAL S3576 : STD_LOGIC;
    SIGNAL S3577 : STD_LOGIC;
    SIGNAL S3578 : STD_LOGIC;
    SIGNAL S3579 : STD_LOGIC;
    SIGNAL S3580 : STD_LOGIC;
    SIGNAL S3581 : STD_LOGIC;
    SIGNAL S3582 : STD_LOGIC;
    SIGNAL S3583 : STD_LOGIC;
    SIGNAL S3584 : STD_LOGIC;
    SIGNAL S3585 : STD_LOGIC;
    SIGNAL S3586 : STD_LOGIC;
    SIGNAL S3587 : STD_LOGIC;
    SIGNAL S3588 : STD_LOGIC;
    SIGNAL S3589 : STD_LOGIC;
    SIGNAL S3590 : STD_LOGIC;
    SIGNAL S3591 : STD_LOGIC;
    SIGNAL S3592 : STD_LOGIC;
    SIGNAL S3593 : STD_LOGIC;
    SIGNAL S3594 : STD_LOGIC;
    SIGNAL S3595 : STD_LOGIC;
    SIGNAL S3596 : STD_LOGIC;
    SIGNAL S3597 : STD_LOGIC;
    SIGNAL S3598 : STD_LOGIC;
    SIGNAL S3599 : STD_LOGIC;
    SIGNAL S3600 : STD_LOGIC;
    SIGNAL S3601 : STD_LOGIC;
    SIGNAL S3602 : STD_LOGIC;
    SIGNAL S3603 : STD_LOGIC;
    SIGNAL S3604 : STD_LOGIC;
    SIGNAL S3605 : STD_LOGIC;
    SIGNAL S3606 : STD_LOGIC;
    SIGNAL S3607 : STD_LOGIC;
    SIGNAL S3608 : STD_LOGIC;
    SIGNAL S3609 : STD_LOGIC;
    SIGNAL S3610 : STD_LOGIC;
    SIGNAL S3611 : STD_LOGIC;
    SIGNAL S3612 : STD_LOGIC;
    SIGNAL S3613 : STD_LOGIC;
    SIGNAL S3614 : STD_LOGIC;
    SIGNAL S3615 : STD_LOGIC;
    SIGNAL S3616 : STD_LOGIC;
    SIGNAL S3617 : STD_LOGIC;
    SIGNAL S3618 : STD_LOGIC;
    SIGNAL S3619 : STD_LOGIC;
    SIGNAL S3620 : STD_LOGIC;
    SIGNAL S3621 : STD_LOGIC;
    SIGNAL S3622 : STD_LOGIC;
    SIGNAL S3623 : STD_LOGIC;
    SIGNAL S3624 : STD_LOGIC;
    SIGNAL S3625 : STD_LOGIC;
    SIGNAL S3626 : STD_LOGIC;
    SIGNAL S3627 : STD_LOGIC;
    SIGNAL S3628 : STD_LOGIC;
    SIGNAL S3629 : STD_LOGIC;
    SIGNAL S3630 : STD_LOGIC;
    SIGNAL S3631 : STD_LOGIC;
    SIGNAL S3632 : STD_LOGIC;
    SIGNAL S3633 : STD_LOGIC;
    SIGNAL S3634 : STD_LOGIC;
    SIGNAL S3635 : STD_LOGIC;
    SIGNAL S3636 : STD_LOGIC;
    SIGNAL S3637 : STD_LOGIC;
    SIGNAL S3638 : STD_LOGIC;
    SIGNAL S3639 : STD_LOGIC;
    SIGNAL S3640 : STD_LOGIC;
    SIGNAL S3641 : STD_LOGIC;
    SIGNAL S3642 : STD_LOGIC;
    SIGNAL S3643 : STD_LOGIC;
    SIGNAL S3644 : STD_LOGIC;
    SIGNAL S3645 : STD_LOGIC;
    SIGNAL S3646 : STD_LOGIC;
    SIGNAL S3647 : STD_LOGIC;
    SIGNAL S3648 : STD_LOGIC;
    SIGNAL S3649 : STD_LOGIC;
    SIGNAL S3650 : STD_LOGIC;
    SIGNAL S3651 : STD_LOGIC;
    SIGNAL S3652 : STD_LOGIC;
    SIGNAL S3653 : STD_LOGIC;
    SIGNAL S3654 : STD_LOGIC;
    SIGNAL S3655 : STD_LOGIC;
    SIGNAL S3656 : STD_LOGIC;
    SIGNAL S3657 : STD_LOGIC;
    SIGNAL S3658 : STD_LOGIC;
    SIGNAL S3659 : STD_LOGIC;
    SIGNAL S3660 : STD_LOGIC;
    SIGNAL S3661 : STD_LOGIC;
    SIGNAL S3662 : STD_LOGIC;
    SIGNAL S3663 : STD_LOGIC;
    SIGNAL S3664 : STD_LOGIC;
    SIGNAL S3665 : STD_LOGIC;
    SIGNAL S3666 : STD_LOGIC;
    SIGNAL S3667 : STD_LOGIC;
    SIGNAL S3668 : STD_LOGIC;
    SIGNAL S3669 : STD_LOGIC;
    SIGNAL S3670 : STD_LOGIC;
    SIGNAL S3671 : STD_LOGIC;
    SIGNAL S3672 : STD_LOGIC;
    SIGNAL S3673 : STD_LOGIC;
    SIGNAL S3674 : STD_LOGIC;
    SIGNAL S3675 : STD_LOGIC;
    SIGNAL S3676 : STD_LOGIC;
    SIGNAL S3677 : STD_LOGIC;
    SIGNAL S3678 : STD_LOGIC;
    SIGNAL S3679 : STD_LOGIC;
    SIGNAL S3680 : STD_LOGIC;
    SIGNAL S3681 : STD_LOGIC;
    SIGNAL S3682 : STD_LOGIC;
    SIGNAL S3683 : STD_LOGIC;
    SIGNAL S3684 : STD_LOGIC;
    SIGNAL S3685 : STD_LOGIC;
    SIGNAL S3686 : STD_LOGIC;
    SIGNAL S3687 : STD_LOGIC;
    SIGNAL S3688 : STD_LOGIC;
    SIGNAL S3689 : STD_LOGIC;
    SIGNAL S3690 : STD_LOGIC;
    SIGNAL S3691 : STD_LOGIC;
    SIGNAL S3692 : STD_LOGIC;
    SIGNAL S3693 : STD_LOGIC;
    SIGNAL S3694 : STD_LOGIC;
    SIGNAL S3695 : STD_LOGIC;
    SIGNAL S3696 : STD_LOGIC;
    SIGNAL S3697 : STD_LOGIC;
    SIGNAL S3698 : STD_LOGIC;
    SIGNAL S3699 : STD_LOGIC;
    SIGNAL S3700 : STD_LOGIC;
    SIGNAL S3701 : STD_LOGIC;
    SIGNAL S3702 : STD_LOGIC;
    SIGNAL S3703 : STD_LOGIC;
    SIGNAL S3704 : STD_LOGIC;
    SIGNAL S3705 : STD_LOGIC;
    SIGNAL S3706 : STD_LOGIC;
    SIGNAL S3707 : STD_LOGIC;
    SIGNAL S3708 : STD_LOGIC;
    SIGNAL S3709 : STD_LOGIC;
    SIGNAL S3710 : STD_LOGIC;
    SIGNAL S3711 : STD_LOGIC;
    SIGNAL S3712 : STD_LOGIC;
    SIGNAL S3713 : STD_LOGIC;
    SIGNAL S3714 : STD_LOGIC;
    SIGNAL S3715 : STD_LOGIC;
    SIGNAL S3716 : STD_LOGIC;
    SIGNAL S3717 : STD_LOGIC;
    SIGNAL S3718 : STD_LOGIC;
    SIGNAL S3719 : STD_LOGIC;
    SIGNAL S3720 : STD_LOGIC;
    SIGNAL S3721 : STD_LOGIC;
    SIGNAL S3722 : STD_LOGIC;
    SIGNAL S3723 : STD_LOGIC;
    SIGNAL S3724 : STD_LOGIC;
    SIGNAL S3725 : STD_LOGIC;
    SIGNAL S3726 : STD_LOGIC;
    SIGNAL S3727 : STD_LOGIC;
    SIGNAL S3728 : STD_LOGIC;
    SIGNAL S3729 : STD_LOGIC;
    SIGNAL S3730 : STD_LOGIC;
    SIGNAL S3731 : STD_LOGIC;
    SIGNAL S3732 : STD_LOGIC;
    SIGNAL S3733 : STD_LOGIC;
    SIGNAL S3734 : STD_LOGIC;
    SIGNAL S3735 : STD_LOGIC;
    SIGNAL S3736 : STD_LOGIC;
    SIGNAL S3737 : STD_LOGIC;
    SIGNAL S3738 : STD_LOGIC;
    SIGNAL S3739 : STD_LOGIC;
    SIGNAL S3740 : STD_LOGIC;
    SIGNAL S3741 : STD_LOGIC;
    SIGNAL S3742 : STD_LOGIC;
    SIGNAL S3743 : STD_LOGIC;
    SIGNAL S3744 : STD_LOGIC;
    SIGNAL S3745 : STD_LOGIC;
    SIGNAL S3746 : STD_LOGIC;
    SIGNAL S3747 : STD_LOGIC;
    SIGNAL S3748 : STD_LOGIC;
    SIGNAL S3749 : STD_LOGIC;
    SIGNAL S3750 : STD_LOGIC;
    SIGNAL S3751 : STD_LOGIC;
    SIGNAL S3752 : STD_LOGIC;
    SIGNAL S3753 : STD_LOGIC;
    SIGNAL S3754 : STD_LOGIC;
    SIGNAL S3755 : STD_LOGIC;
    SIGNAL S3756 : STD_LOGIC;
    SIGNAL S3757 : STD_LOGIC;
    SIGNAL S3758 : STD_LOGIC;
    SIGNAL S3759 : STD_LOGIC;
    SIGNAL S3760 : STD_LOGIC;
    SIGNAL S3761 : STD_LOGIC;
    SIGNAL S3762 : STD_LOGIC;
    SIGNAL S3763 : STD_LOGIC;
    SIGNAL S3764 : STD_LOGIC;
    SIGNAL S3765 : STD_LOGIC;
    SIGNAL S3766 : STD_LOGIC;
    SIGNAL S3767 : STD_LOGIC;
    SIGNAL S3768 : STD_LOGIC;
    SIGNAL S3769 : STD_LOGIC;
    SIGNAL S3770 : STD_LOGIC;
    SIGNAL S3771 : STD_LOGIC;
    SIGNAL S3772 : STD_LOGIC;
    SIGNAL S3773 : STD_LOGIC;
    SIGNAL S3774 : STD_LOGIC;
    SIGNAL S3775 : STD_LOGIC;
    SIGNAL S3776 : STD_LOGIC;
    SIGNAL S3777 : STD_LOGIC;
    SIGNAL S3778 : STD_LOGIC;
    SIGNAL S3779 : STD_LOGIC;
    SIGNAL S3780 : STD_LOGIC;
    SIGNAL S3781 : STD_LOGIC;
    SIGNAL S3782 : STD_LOGIC;
    SIGNAL S3783 : STD_LOGIC;
    SIGNAL S3784 : STD_LOGIC;
    SIGNAL S3785 : STD_LOGIC;
    SIGNAL S3786 : STD_LOGIC;
    SIGNAL S3787 : STD_LOGIC;
    SIGNAL S3788 : STD_LOGIC;
    SIGNAL S3789 : STD_LOGIC;
    SIGNAL S3790 : STD_LOGIC;
    SIGNAL S3791 : STD_LOGIC;
    SIGNAL S3792 : STD_LOGIC;
    SIGNAL S3793 : STD_LOGIC;
    SIGNAL S3794 : STD_LOGIC;
    SIGNAL S3795 : STD_LOGIC;
    SIGNAL S3796 : STD_LOGIC;
    SIGNAL S3797 : STD_LOGIC;
    SIGNAL S3798 : STD_LOGIC;
    SIGNAL S3799 : STD_LOGIC;
    SIGNAL S3800 : STD_LOGIC;
    SIGNAL S3801 : STD_LOGIC;
    SIGNAL S3802 : STD_LOGIC;
    SIGNAL S3803 : STD_LOGIC;
    SIGNAL S3804 : STD_LOGIC;
    SIGNAL S3805 : STD_LOGIC;
    SIGNAL S3806 : STD_LOGIC;
    SIGNAL S3807 : STD_LOGIC;
    SIGNAL S3808 : STD_LOGIC;
    SIGNAL S3809 : STD_LOGIC;
    SIGNAL S3810 : STD_LOGIC;
    SIGNAL S3811 : STD_LOGIC;
    SIGNAL S3812 : STD_LOGIC;
    SIGNAL S3813 : STD_LOGIC;
    SIGNAL S3814 : STD_LOGIC;
    SIGNAL S3815 : STD_LOGIC;
    SIGNAL S3816 : STD_LOGIC;
    SIGNAL S3817 : STD_LOGIC;
    SIGNAL S3818 : STD_LOGIC;
    SIGNAL S3819 : STD_LOGIC;
    SIGNAL S3820 : STD_LOGIC;
    SIGNAL S3821 : STD_LOGIC;
    SIGNAL S3822 : STD_LOGIC;
    SIGNAL S3823 : STD_LOGIC;
    SIGNAL S3824 : STD_LOGIC;
    SIGNAL S3825 : STD_LOGIC;
    SIGNAL S3826 : STD_LOGIC;
    SIGNAL S3827 : STD_LOGIC;
    SIGNAL S3828 : STD_LOGIC;
    SIGNAL S3829 : STD_LOGIC;
    SIGNAL S3830 : STD_LOGIC;
    SIGNAL S3831 : STD_LOGIC;
    SIGNAL S3832 : STD_LOGIC;
    SIGNAL S3833 : STD_LOGIC;
    SIGNAL S3834 : STD_LOGIC;
    SIGNAL S3835 : STD_LOGIC;
    SIGNAL S3836 : STD_LOGIC;
    SIGNAL S3837 : STD_LOGIC;
    SIGNAL S3838 : STD_LOGIC;
    SIGNAL S3839 : STD_LOGIC;
    SIGNAL S3840 : STD_LOGIC;
    SIGNAL S3841 : STD_LOGIC;
    SIGNAL S3842 : STD_LOGIC;
    SIGNAL S3843 : STD_LOGIC;
    SIGNAL S3844 : STD_LOGIC;
    SIGNAL S3845 : STD_LOGIC;
    SIGNAL S3846 : STD_LOGIC;
    SIGNAL S3847 : STD_LOGIC;
    SIGNAL S3848 : STD_LOGIC;
    SIGNAL S3849 : STD_LOGIC;
    SIGNAL S3850 : STD_LOGIC;
    SIGNAL S3851 : STD_LOGIC;
    SIGNAL S3852 : STD_LOGIC;
    SIGNAL S3853 : STD_LOGIC;
    SIGNAL S3854 : STD_LOGIC;
    SIGNAL S3855 : STD_LOGIC;
    SIGNAL S3856 : STD_LOGIC;
    SIGNAL S3857 : STD_LOGIC;
    SIGNAL S3858 : STD_LOGIC;
    SIGNAL S3859 : STD_LOGIC;
    SIGNAL S3860 : STD_LOGIC;
    SIGNAL S3861 : STD_LOGIC;
    SIGNAL S3862 : STD_LOGIC;
    SIGNAL S3863 : STD_LOGIC;
    SIGNAL S3864 : STD_LOGIC;
    SIGNAL S3865 : STD_LOGIC;
    SIGNAL S3866 : STD_LOGIC;
    SIGNAL S3867 : STD_LOGIC;
    SIGNAL S3868 : STD_LOGIC;
    SIGNAL S3869 : STD_LOGIC;
    SIGNAL S3870 : STD_LOGIC;
    SIGNAL S3871 : STD_LOGIC;
    SIGNAL S3872 : STD_LOGIC;
    SIGNAL S3873 : STD_LOGIC;
    SIGNAL S3874 : STD_LOGIC;
    SIGNAL S3875 : STD_LOGIC;
    SIGNAL S3876 : STD_LOGIC;
    SIGNAL S3877 : STD_LOGIC;
    SIGNAL S3878 : STD_LOGIC;
    SIGNAL S3879 : STD_LOGIC;
    SIGNAL S3880 : STD_LOGIC;
    SIGNAL S3881 : STD_LOGIC;
    SIGNAL S3882 : STD_LOGIC;
    SIGNAL S3883 : STD_LOGIC;
    SIGNAL S3884 : STD_LOGIC;
    SIGNAL S3885 : STD_LOGIC;
    SIGNAL S3886 : STD_LOGIC;
    SIGNAL S3887 : STD_LOGIC;
    SIGNAL S3888 : STD_LOGIC;
    SIGNAL S3889 : STD_LOGIC;
    SIGNAL S3890 : STD_LOGIC;
    SIGNAL S3891 : STD_LOGIC;
    SIGNAL S3892 : STD_LOGIC;
    SIGNAL S3893 : STD_LOGIC;
    SIGNAL S3894 : STD_LOGIC;
    SIGNAL S3895 : STD_LOGIC;
    SIGNAL S3896 : STD_LOGIC;
    SIGNAL S3897 : STD_LOGIC;
    SIGNAL S3898 : STD_LOGIC;
    SIGNAL S3899 : STD_LOGIC;
    SIGNAL S3900 : STD_LOGIC;
    SIGNAL S3901 : STD_LOGIC;
    SIGNAL S3902 : STD_LOGIC;
    SIGNAL S3903 : STD_LOGIC;
    SIGNAL S3904 : STD_LOGIC;
    SIGNAL S3905 : STD_LOGIC;
    SIGNAL S3906 : STD_LOGIC;
    SIGNAL S3907 : STD_LOGIC;
    SIGNAL S3908 : STD_LOGIC;
    SIGNAL S3909 : STD_LOGIC;
    SIGNAL S3910 : STD_LOGIC;
    SIGNAL S3911 : STD_LOGIC;
    SIGNAL S3912 : STD_LOGIC;
    SIGNAL S3913 : STD_LOGIC;
    SIGNAL S3914 : STD_LOGIC;
    SIGNAL S3915 : STD_LOGIC;
    SIGNAL S3916 : STD_LOGIC;
    SIGNAL S3917 : STD_LOGIC;
    SIGNAL S3918 : STD_LOGIC;
    SIGNAL S3919 : STD_LOGIC;
    SIGNAL S3920 : STD_LOGIC;
    SIGNAL S3921 : STD_LOGIC;
    SIGNAL S3922 : STD_LOGIC;
    SIGNAL S3923 : STD_LOGIC;
    SIGNAL S3924 : STD_LOGIC;
    SIGNAL S3925 : STD_LOGIC;
    SIGNAL S3926 : STD_LOGIC;
    SIGNAL S3927 : STD_LOGIC;
    SIGNAL S3928 : STD_LOGIC;
    SIGNAL S3929 : STD_LOGIC;
    SIGNAL S3930 : STD_LOGIC;
    SIGNAL S3931 : STD_LOGIC;
    SIGNAL S3932 : STD_LOGIC;
    SIGNAL S3933 : STD_LOGIC;
    SIGNAL S3934 : STD_LOGIC;
    SIGNAL S3935 : STD_LOGIC;
    SIGNAL S3936 : STD_LOGIC;
    SIGNAL S3937 : STD_LOGIC;
    SIGNAL S3938 : STD_LOGIC;
    SIGNAL S3939 : STD_LOGIC;
    SIGNAL S3940 : STD_LOGIC;
    SIGNAL S3941 : STD_LOGIC;
    SIGNAL S3942 : STD_LOGIC;
    SIGNAL S3943 : STD_LOGIC;
    SIGNAL S3944 : STD_LOGIC;
    SIGNAL S3945 : STD_LOGIC;
    SIGNAL S3946 : STD_LOGIC;
    SIGNAL S3947 : STD_LOGIC;
    SIGNAL S3948 : STD_LOGIC;
    SIGNAL S3949 : STD_LOGIC;
    SIGNAL S3950 : STD_LOGIC;
    SIGNAL S3951 : STD_LOGIC;
    SIGNAL S3952 : STD_LOGIC;
    SIGNAL S3953 : STD_LOGIC;
    SIGNAL S3954 : STD_LOGIC;
    SIGNAL S3955 : STD_LOGIC;
    SIGNAL S3956 : STD_LOGIC;
    SIGNAL S3957 : STD_LOGIC;
    SIGNAL S3958 : STD_LOGIC;
    SIGNAL S3959 : STD_LOGIC;
    SIGNAL S3960 : STD_LOGIC;
    SIGNAL S3961 : STD_LOGIC;
    SIGNAL S3962 : STD_LOGIC;
    SIGNAL S3963 : STD_LOGIC;
    SIGNAL S3964 : STD_LOGIC;
    SIGNAL S3965 : STD_LOGIC;
    SIGNAL S3966 : STD_LOGIC;
    SIGNAL S3967 : STD_LOGIC;
    SIGNAL S3968 : STD_LOGIC;
    SIGNAL S3969 : STD_LOGIC;
    SIGNAL S3970 : STD_LOGIC;
    SIGNAL S3971 : STD_LOGIC;
    SIGNAL S3972 : STD_LOGIC;
    SIGNAL S3973 : STD_LOGIC;
    SIGNAL S3974 : STD_LOGIC;
    SIGNAL S3975 : STD_LOGIC;
    SIGNAL S3976 : STD_LOGIC;
    SIGNAL S3977 : STD_LOGIC;
    SIGNAL S3978 : STD_LOGIC;
    SIGNAL S3979 : STD_LOGIC;
    SIGNAL S3980 : STD_LOGIC;
    SIGNAL S3981 : STD_LOGIC;
    SIGNAL S3982 : STD_LOGIC;
    SIGNAL S3983 : STD_LOGIC;
    SIGNAL S3984 : STD_LOGIC;
    SIGNAL S3985 : STD_LOGIC;
    SIGNAL S3986 : STD_LOGIC;
    SIGNAL S3987 : STD_LOGIC;
    SIGNAL S3988 : STD_LOGIC;
    SIGNAL S3989 : STD_LOGIC;
    SIGNAL S3990 : STD_LOGIC;
    SIGNAL S3991 : STD_LOGIC;
    SIGNAL S3992 : STD_LOGIC;
    SIGNAL S3993 : STD_LOGIC;
    SIGNAL S3994 : STD_LOGIC;
    SIGNAL S3995 : STD_LOGIC;
    SIGNAL S3996 : STD_LOGIC;
    SIGNAL S3997 : STD_LOGIC;
    SIGNAL S3998 : STD_LOGIC;
    SIGNAL S3999 : STD_LOGIC;
    SIGNAL S4000 : STD_LOGIC;
    SIGNAL S4001 : STD_LOGIC;
    SIGNAL S4002 : STD_LOGIC;
    SIGNAL S4003 : STD_LOGIC;
    SIGNAL S4004 : STD_LOGIC;
    SIGNAL S4005 : STD_LOGIC;
    SIGNAL S4006 : STD_LOGIC;
    SIGNAL S4007 : STD_LOGIC;
    SIGNAL S4008 : STD_LOGIC;
    SIGNAL S4009 : STD_LOGIC;
    SIGNAL S4010 : STD_LOGIC;
    SIGNAL S4011 : STD_LOGIC;
    SIGNAL S4012 : STD_LOGIC;
    SIGNAL S4013 : STD_LOGIC;
    SIGNAL S4014 : STD_LOGIC;
    SIGNAL S4015 : STD_LOGIC;
    SIGNAL S4016 : STD_LOGIC;
    SIGNAL S4017 : STD_LOGIC;
    SIGNAL S4018 : STD_LOGIC;
    SIGNAL S4019 : STD_LOGIC;
    SIGNAL S4020 : STD_LOGIC;
    SIGNAL S4021 : STD_LOGIC;
    SIGNAL S4022 : STD_LOGIC;
    SIGNAL S4023 : STD_LOGIC;
    SIGNAL S4024 : STD_LOGIC;
    SIGNAL S4025 : STD_LOGIC;
    SIGNAL S4026 : STD_LOGIC;
    SIGNAL S4027 : STD_LOGIC;
    SIGNAL S4028 : STD_LOGIC;
    SIGNAL S4029 : STD_LOGIC;
    SIGNAL S4030 : STD_LOGIC;
    SIGNAL S4031 : STD_LOGIC;
    SIGNAL S4032 : STD_LOGIC;
    SIGNAL S4033 : STD_LOGIC;
    SIGNAL S4034 : STD_LOGIC;
    SIGNAL S4035 : STD_LOGIC;
    SIGNAL S4036 : STD_LOGIC;
    SIGNAL S4037 : STD_LOGIC;
    SIGNAL S4038 : STD_LOGIC;
    SIGNAL S4039 : STD_LOGIC;
    SIGNAL S4040 : STD_LOGIC;
    SIGNAL S4041 : STD_LOGIC;
    SIGNAL S4042 : STD_LOGIC;
    SIGNAL S4043 : STD_LOGIC;
    SIGNAL S4044 : STD_LOGIC;
    SIGNAL S4045 : STD_LOGIC;
    SIGNAL S4046 : STD_LOGIC;
    SIGNAL S4047 : STD_LOGIC;
    SIGNAL S4048 : STD_LOGIC;
    SIGNAL S4049 : STD_LOGIC;
    SIGNAL S4050 : STD_LOGIC;
    SIGNAL S4051 : STD_LOGIC;
    SIGNAL S4052 : STD_LOGIC;
    SIGNAL S4053 : STD_LOGIC;
    SIGNAL S4054 : STD_LOGIC;
    SIGNAL S4055 : STD_LOGIC;
    SIGNAL S4056 : STD_LOGIC;
    SIGNAL S4057 : STD_LOGIC;
    SIGNAL S4058 : STD_LOGIC;
    SIGNAL S4059 : STD_LOGIC;
    SIGNAL S4060 : STD_LOGIC;
    SIGNAL S4061 : STD_LOGIC;
    SIGNAL S4062 : STD_LOGIC;
    SIGNAL S4063 : STD_LOGIC;
    SIGNAL S4064 : STD_LOGIC;
    SIGNAL S4065 : STD_LOGIC;
    SIGNAL S4066 : STD_LOGIC;
    SIGNAL S4067 : STD_LOGIC;
    SIGNAL S4068 : STD_LOGIC;
    SIGNAL S4069 : STD_LOGIC;
    SIGNAL S4070 : STD_LOGIC;
    SIGNAL S4071 : STD_LOGIC;
    SIGNAL S4072 : STD_LOGIC;
    SIGNAL S4073 : STD_LOGIC;
    SIGNAL S4074 : STD_LOGIC;
    SIGNAL S4075 : STD_LOGIC;
    SIGNAL S4076 : STD_LOGIC;
    SIGNAL S4077 : STD_LOGIC;
    SIGNAL S4078 : STD_LOGIC;
    SIGNAL S4079 : STD_LOGIC;
    SIGNAL S4080 : STD_LOGIC;
    SIGNAL S4081 : STD_LOGIC;
    SIGNAL S4082 : STD_LOGIC;
    SIGNAL S4083 : STD_LOGIC;
    SIGNAL S4084 : STD_LOGIC;
    SIGNAL S4085 : STD_LOGIC;
    SIGNAL S4086 : STD_LOGIC;
    SIGNAL S4087 : STD_LOGIC;
    SIGNAL S4088 : STD_LOGIC;
    SIGNAL S4089 : STD_LOGIC;
    SIGNAL S4090 : STD_LOGIC;
    SIGNAL S4091 : STD_LOGIC;
    SIGNAL S4092 : STD_LOGIC;
    SIGNAL S4093 : STD_LOGIC;
    SIGNAL S4094 : STD_LOGIC;
    SIGNAL S4095 : STD_LOGIC;
    SIGNAL S4096 : STD_LOGIC;
    SIGNAL S4097 : STD_LOGIC;
    SIGNAL S4098 : STD_LOGIC;
    SIGNAL S4099 : STD_LOGIC;
    SIGNAL S4100 : STD_LOGIC;
    SIGNAL S4101 : STD_LOGIC;
    SIGNAL S4102 : STD_LOGIC;
    SIGNAL S4103 : STD_LOGIC;
    SIGNAL S4104 : STD_LOGIC;
    SIGNAL S4105 : STD_LOGIC;
    SIGNAL S4106 : STD_LOGIC;
    SIGNAL S4107 : STD_LOGIC;
    SIGNAL S4108 : STD_LOGIC;
    SIGNAL S4109 : STD_LOGIC;
    SIGNAL S4110 : STD_LOGIC;
    SIGNAL S4111 : STD_LOGIC;
    SIGNAL S4112 : STD_LOGIC;
    SIGNAL S4113 : STD_LOGIC;
    SIGNAL S4114 : STD_LOGIC;
    SIGNAL S4115 : STD_LOGIC;
    SIGNAL S4116 : STD_LOGIC;
    SIGNAL S4117 : STD_LOGIC;
    SIGNAL S4118 : STD_LOGIC;
    SIGNAL S4119 : STD_LOGIC;
    SIGNAL S4120 : STD_LOGIC;
    SIGNAL S4121 : STD_LOGIC;
    SIGNAL S4122 : STD_LOGIC;
    SIGNAL S4123 : STD_LOGIC;
    SIGNAL S4124 : STD_LOGIC;
    SIGNAL S4125 : STD_LOGIC;
    SIGNAL S4126 : STD_LOGIC;
    SIGNAL S4127 : STD_LOGIC;
    SIGNAL S4128 : STD_LOGIC;
    SIGNAL S4129 : STD_LOGIC;
    SIGNAL S4130 : STD_LOGIC;
    SIGNAL S4131 : STD_LOGIC;
    SIGNAL S4132 : STD_LOGIC;
    SIGNAL S4133 : STD_LOGIC;
    SIGNAL S4134 : STD_LOGIC;
    SIGNAL S4135 : STD_LOGIC;
    SIGNAL S4136 : STD_LOGIC;
    SIGNAL S4137 : STD_LOGIC;
    SIGNAL S4138 : STD_LOGIC;
    SIGNAL S4139 : STD_LOGIC;
    SIGNAL S4140 : STD_LOGIC;
    SIGNAL S4141 : STD_LOGIC;
    SIGNAL S4142 : STD_LOGIC;
    SIGNAL S4143 : STD_LOGIC;
    SIGNAL S4144 : STD_LOGIC;
    SIGNAL S4145 : STD_LOGIC;
    SIGNAL S4146 : STD_LOGIC;
    SIGNAL S4147 : STD_LOGIC;
    SIGNAL S4148 : STD_LOGIC;
    SIGNAL S4149 : STD_LOGIC;
    SIGNAL S4150 : STD_LOGIC;
    SIGNAL S4151 : STD_LOGIC;
    SIGNAL S4152 : STD_LOGIC;
    SIGNAL S4153 : STD_LOGIC;
    SIGNAL S4154 : STD_LOGIC;
    SIGNAL S4155 : STD_LOGIC;
    SIGNAL S4156 : STD_LOGIC;
    SIGNAL S4157 : STD_LOGIC;
    SIGNAL S4158 : STD_LOGIC;
    SIGNAL S4159 : STD_LOGIC;
    SIGNAL S4160 : STD_LOGIC;
    SIGNAL S4161 : STD_LOGIC;
    SIGNAL S4162 : STD_LOGIC;
    SIGNAL S4163 : STD_LOGIC;
    SIGNAL S4164 : STD_LOGIC;
    SIGNAL S4165 : STD_LOGIC;
    SIGNAL S4166 : STD_LOGIC;
    SIGNAL S4167 : STD_LOGIC;
    SIGNAL S4168 : STD_LOGIC;
    SIGNAL S4169 : STD_LOGIC;
    SIGNAL S4170 : STD_LOGIC;
    SIGNAL S4171 : STD_LOGIC;
    SIGNAL S4172 : STD_LOGIC;
    SIGNAL S4173 : STD_LOGIC;
    SIGNAL S4174 : STD_LOGIC;
    SIGNAL S4175 : STD_LOGIC;
    SIGNAL S4176 : STD_LOGIC;
    SIGNAL S4177 : STD_LOGIC;
    SIGNAL S4178 : STD_LOGIC;
    SIGNAL S4179 : STD_LOGIC;
    SIGNAL S4180 : STD_LOGIC;
    SIGNAL S4181 : STD_LOGIC;
    SIGNAL S4182 : STD_LOGIC;
    SIGNAL S4183 : STD_LOGIC;
    SIGNAL S4184 : STD_LOGIC;
    SIGNAL S4185 : STD_LOGIC;
    SIGNAL S4186 : STD_LOGIC;
    SIGNAL S4187 : STD_LOGIC;
    SIGNAL S4188 : STD_LOGIC;
    SIGNAL S4189 : STD_LOGIC;
    SIGNAL S4190 : STD_LOGIC;
    SIGNAL S4191 : STD_LOGIC;
    SIGNAL S4192 : STD_LOGIC;
    SIGNAL S4193 : STD_LOGIC;
    SIGNAL S4194 : STD_LOGIC;
    SIGNAL S4195 : STD_LOGIC;
    SIGNAL S4196 : STD_LOGIC;
    SIGNAL S4197 : STD_LOGIC;
    SIGNAL S4198 : STD_LOGIC;
    SIGNAL S4199 : STD_LOGIC;
    SIGNAL S4200 : STD_LOGIC;
    SIGNAL S4201 : STD_LOGIC;
    SIGNAL S4202 : STD_LOGIC;
    SIGNAL S4203 : STD_LOGIC;
    SIGNAL S4204 : STD_LOGIC;
    SIGNAL S4205 : STD_LOGIC;
    SIGNAL S4206 : STD_LOGIC;
    SIGNAL S4207 : STD_LOGIC;
    SIGNAL S4208 : STD_LOGIC;
    SIGNAL S4209 : STD_LOGIC;
    SIGNAL S4210 : STD_LOGIC;
    SIGNAL S4211 : STD_LOGIC;
    SIGNAL S4212 : STD_LOGIC;
    SIGNAL S4213 : STD_LOGIC;
    SIGNAL S4214 : STD_LOGIC;
    SIGNAL S4215 : STD_LOGIC;
    SIGNAL S4216 : STD_LOGIC;
    SIGNAL S4217 : STD_LOGIC;
    SIGNAL S4218 : STD_LOGIC;
    SIGNAL S4219 : STD_LOGIC;
    SIGNAL S4220 : STD_LOGIC;
    SIGNAL S4221 : STD_LOGIC;
    SIGNAL S4222 : STD_LOGIC;
    SIGNAL S4223 : STD_LOGIC;
    SIGNAL S4224 : STD_LOGIC;
    SIGNAL S4225 : STD_LOGIC;
    SIGNAL S4226 : STD_LOGIC;
    SIGNAL S4227 : STD_LOGIC;
    SIGNAL S4228 : STD_LOGIC;
    SIGNAL S4229 : STD_LOGIC;
    SIGNAL S4230 : STD_LOGIC;
    SIGNAL S4231 : STD_LOGIC;
    SIGNAL S4232 : STD_LOGIC;
    SIGNAL S4233 : STD_LOGIC;
    SIGNAL S4234 : STD_LOGIC;
    SIGNAL S4235 : STD_LOGIC;
    SIGNAL S4236 : STD_LOGIC;
    SIGNAL S4237 : STD_LOGIC;
    SIGNAL S4238 : STD_LOGIC;
    SIGNAL S4239 : STD_LOGIC;
    SIGNAL S4240 : STD_LOGIC;
    SIGNAL S4241 : STD_LOGIC;
    SIGNAL S4242 : STD_LOGIC;
    SIGNAL S4243 : STD_LOGIC;
    SIGNAL S4244 : STD_LOGIC;
    SIGNAL S4245 : STD_LOGIC;
    SIGNAL S4246 : STD_LOGIC;
    SIGNAL S4247 : STD_LOGIC;
    SIGNAL S4248 : STD_LOGIC;
    SIGNAL S4249 : STD_LOGIC;
    SIGNAL S4250 : STD_LOGIC;
    SIGNAL S4251 : STD_LOGIC;
    SIGNAL S4252 : STD_LOGIC;
    SIGNAL S4253 : STD_LOGIC;
    SIGNAL S4254 : STD_LOGIC;
    SIGNAL S4255 : STD_LOGIC;
    SIGNAL S4256 : STD_LOGIC;
    SIGNAL S4257 : STD_LOGIC;
    SIGNAL S4258 : STD_LOGIC;
    SIGNAL S4259 : STD_LOGIC;
    SIGNAL S4260 : STD_LOGIC;
    SIGNAL S4261 : STD_LOGIC;
    SIGNAL S4262 : STD_LOGIC;
    SIGNAL S4263 : STD_LOGIC;
    SIGNAL S4264 : STD_LOGIC;
    SIGNAL S4265 : STD_LOGIC;
    SIGNAL S4266 : STD_LOGIC;
    SIGNAL S4267 : STD_LOGIC;
    SIGNAL S4268 : STD_LOGIC;
    SIGNAL S4269 : STD_LOGIC;
    SIGNAL S4270 : STD_LOGIC;
    SIGNAL S4271 : STD_LOGIC;
    SIGNAL S4272 : STD_LOGIC;
    SIGNAL S4273 : STD_LOGIC;
    SIGNAL S4274 : STD_LOGIC;
    SIGNAL S4275 : STD_LOGIC;
    SIGNAL S4276 : STD_LOGIC;
    SIGNAL S4277 : STD_LOGIC;
    SIGNAL S4278 : STD_LOGIC;
    SIGNAL S4279 : STD_LOGIC;
    SIGNAL S4280 : STD_LOGIC;
    SIGNAL S4281 : STD_LOGIC;
    SIGNAL S4282 : STD_LOGIC;
    SIGNAL S4283 : STD_LOGIC;
    SIGNAL S4284 : STD_LOGIC;
    SIGNAL S4285 : STD_LOGIC;
    SIGNAL S4286 : STD_LOGIC;
    SIGNAL S4287 : STD_LOGIC;
    SIGNAL S4288 : STD_LOGIC;
    SIGNAL S4289 : STD_LOGIC;
    SIGNAL S4290 : STD_LOGIC;
    SIGNAL S4291 : STD_LOGIC;
    SIGNAL S4292 : STD_LOGIC;
    SIGNAL S4293 : STD_LOGIC;
    SIGNAL S4294 : STD_LOGIC;
    SIGNAL S4295 : STD_LOGIC;
    SIGNAL S4296 : STD_LOGIC;
    SIGNAL S4297 : STD_LOGIC;
    SIGNAL S4298 : STD_LOGIC;
    SIGNAL S4299 : STD_LOGIC;
    SIGNAL S4300 : STD_LOGIC;
    SIGNAL S4301 : STD_LOGIC;
    SIGNAL S4302 : STD_LOGIC;
    SIGNAL S4303 : STD_LOGIC;
    SIGNAL S4304 : STD_LOGIC;
    SIGNAL S4305 : STD_LOGIC;
    SIGNAL S4306 : STD_LOGIC;
    SIGNAL S4307 : STD_LOGIC;
    SIGNAL S4308 : STD_LOGIC;
    SIGNAL S4309 : STD_LOGIC;
    SIGNAL S4310 : STD_LOGIC;
    SIGNAL S4311 : STD_LOGIC;
    SIGNAL S4312 : STD_LOGIC;
    SIGNAL S4313 : STD_LOGIC;
    SIGNAL S4314 : STD_LOGIC;
    SIGNAL S4315 : STD_LOGIC;
    SIGNAL S4316 : STD_LOGIC;
    SIGNAL S4317 : STD_LOGIC;
    SIGNAL S4318 : STD_LOGIC;
    SIGNAL S4319 : STD_LOGIC;
    SIGNAL S4320 : STD_LOGIC;
    SIGNAL S4321 : STD_LOGIC;
    SIGNAL S4322 : STD_LOGIC;
    SIGNAL S4323 : STD_LOGIC;
    SIGNAL S4324 : STD_LOGIC;
    SIGNAL S4325 : STD_LOGIC;
    SIGNAL S4326 : STD_LOGIC;
    SIGNAL S4327 : STD_LOGIC;
    SIGNAL S4328 : STD_LOGIC;
    SIGNAL S4329 : STD_LOGIC;
    SIGNAL S4330 : STD_LOGIC;
    SIGNAL S4331 : STD_LOGIC;
    SIGNAL S4332 : STD_LOGIC;
    SIGNAL S4333 : STD_LOGIC;
    SIGNAL S4334 : STD_LOGIC;
    SIGNAL S4335 : STD_LOGIC;
    SIGNAL S4336 : STD_LOGIC;
    SIGNAL S4337 : STD_LOGIC;
    SIGNAL S4338 : STD_LOGIC;
    SIGNAL S4339 : STD_LOGIC;
    SIGNAL S4340 : STD_LOGIC;
    SIGNAL S4341 : STD_LOGIC;
    SIGNAL S4342 : STD_LOGIC;
    SIGNAL S4343 : STD_LOGIC;
    SIGNAL S4344 : STD_LOGIC;
    SIGNAL S4345 : STD_LOGIC;
    SIGNAL S4346 : STD_LOGIC;
    SIGNAL S4347 : STD_LOGIC;
    SIGNAL S4348 : STD_LOGIC;
    SIGNAL S4349 : STD_LOGIC;
    SIGNAL S4350 : STD_LOGIC;
    SIGNAL S4351 : STD_LOGIC;
    SIGNAL S4352 : STD_LOGIC;
    SIGNAL S4353 : STD_LOGIC;
    SIGNAL S4354 : STD_LOGIC;
    SIGNAL S4355 : STD_LOGIC;
    SIGNAL S4356 : STD_LOGIC;
    SIGNAL S4357 : STD_LOGIC;
    SIGNAL S4358 : STD_LOGIC;
    SIGNAL S4359 : STD_LOGIC;
    SIGNAL S4360 : STD_LOGIC;
    SIGNAL S4361 : STD_LOGIC;
    SIGNAL S4362 : STD_LOGIC;
    SIGNAL S4363 : STD_LOGIC;
    SIGNAL S4364 : STD_LOGIC;
    SIGNAL S4365 : STD_LOGIC;
    SIGNAL S4366 : STD_LOGIC;
    SIGNAL S4367 : STD_LOGIC;
    SIGNAL S4368 : STD_LOGIC;
    SIGNAL S4369 : STD_LOGIC;
    SIGNAL S4370 : STD_LOGIC;
    SIGNAL S4371 : STD_LOGIC;
    SIGNAL S4372 : STD_LOGIC;
    SIGNAL S4373 : STD_LOGIC;
    SIGNAL S4374 : STD_LOGIC;
    SIGNAL S4375 : STD_LOGIC;
    SIGNAL S4376 : STD_LOGIC;
    SIGNAL S4377 : STD_LOGIC;
    SIGNAL S4378 : STD_LOGIC;
    SIGNAL S4379 : STD_LOGIC;
    SIGNAL S4380 : STD_LOGIC;
    SIGNAL S4381 : STD_LOGIC;
    SIGNAL S4382 : STD_LOGIC;
    SIGNAL S4383 : STD_LOGIC;
    SIGNAL S4384 : STD_LOGIC;
    SIGNAL S4385 : STD_LOGIC;
    SIGNAL S4386 : STD_LOGIC;
    SIGNAL S4387 : STD_LOGIC;
    SIGNAL S4388 : STD_LOGIC;
    SIGNAL S4389 : STD_LOGIC;
    SIGNAL S4390 : STD_LOGIC;
    SIGNAL S4391 : STD_LOGIC;
    SIGNAL S4392 : STD_LOGIC;
    SIGNAL S4393 : STD_LOGIC;
    SIGNAL S4394 : STD_LOGIC;
    SIGNAL S4395 : STD_LOGIC;
    SIGNAL S4396 : STD_LOGIC;
    SIGNAL S4397 : STD_LOGIC;
    SIGNAL S4398 : STD_LOGIC;
    SIGNAL S4399 : STD_LOGIC;
    SIGNAL S4400 : STD_LOGIC;
    SIGNAL S4401 : STD_LOGIC;
    SIGNAL S4402 : STD_LOGIC;
    SIGNAL S4403 : STD_LOGIC;
    SIGNAL S4404 : STD_LOGIC;
    SIGNAL S4405 : STD_LOGIC;
    SIGNAL S4406 : STD_LOGIC;
    SIGNAL S4407 : STD_LOGIC;
    SIGNAL S4408 : STD_LOGIC;
    SIGNAL S4409 : STD_LOGIC;
    SIGNAL S4410 : STD_LOGIC;
    SIGNAL S4411 : STD_LOGIC;
    SIGNAL S4412 : STD_LOGIC;
    SIGNAL S4413 : STD_LOGIC;
    SIGNAL S4414 : STD_LOGIC;
    SIGNAL S4415 : STD_LOGIC;
    SIGNAL S4416 : STD_LOGIC;
    SIGNAL S4417 : STD_LOGIC;
    SIGNAL S4418 : STD_LOGIC;
    SIGNAL S4419 : STD_LOGIC;
    SIGNAL S4420 : STD_LOGIC;
    SIGNAL S4421 : STD_LOGIC;
    SIGNAL S4422 : STD_LOGIC;
    SIGNAL S4423 : STD_LOGIC;
    SIGNAL S4424 : STD_LOGIC;
    SIGNAL S4425 : STD_LOGIC;
    SIGNAL S4426 : STD_LOGIC;
    SIGNAL S4427 : STD_LOGIC;
    SIGNAL S4428 : STD_LOGIC;
    SIGNAL S4429 : STD_LOGIC;
    SIGNAL S4430 : STD_LOGIC;
    SIGNAL S4431 : STD_LOGIC;
    SIGNAL S4432 : STD_LOGIC;
    SIGNAL S4433 : STD_LOGIC;
    SIGNAL S4434 : STD_LOGIC;
    SIGNAL S4435 : STD_LOGIC;
    SIGNAL S4436 : STD_LOGIC;
    SIGNAL S4437 : STD_LOGIC;
    SIGNAL S4438 : STD_LOGIC;
    SIGNAL S4439 : STD_LOGIC;
    SIGNAL S4440 : STD_LOGIC;
    SIGNAL S4441 : STD_LOGIC;
    SIGNAL S4442 : STD_LOGIC;
    SIGNAL S4443 : STD_LOGIC;
    SIGNAL S4444 : STD_LOGIC;
    SIGNAL S4445 : STD_LOGIC;
    SIGNAL S4446 : STD_LOGIC;
    SIGNAL S4447 : STD_LOGIC;
    SIGNAL S4448 : STD_LOGIC;
    SIGNAL S4449 : STD_LOGIC;
    SIGNAL S4450 : STD_LOGIC;
    SIGNAL S4451 : STD_LOGIC;
    SIGNAL S4452 : STD_LOGIC;
    SIGNAL S4453 : STD_LOGIC;
    SIGNAL S4454 : STD_LOGIC;
    SIGNAL S4455 : STD_LOGIC;
    SIGNAL S4456 : STD_LOGIC;
    SIGNAL S4457 : STD_LOGIC;
    SIGNAL S4458 : STD_LOGIC;
    SIGNAL S4459 : STD_LOGIC;
    SIGNAL S4460 : STD_LOGIC;
    SIGNAL S4461 : STD_LOGIC;
    SIGNAL S4462 : STD_LOGIC;
    SIGNAL S4463 : STD_LOGIC;
    SIGNAL S4464 : STD_LOGIC;
    SIGNAL S4465 : STD_LOGIC;
    SIGNAL S4466 : STD_LOGIC;
    SIGNAL S4467 : STD_LOGIC;
    SIGNAL S4468 : STD_LOGIC;
    SIGNAL S4469 : STD_LOGIC;
    SIGNAL S4470 : STD_LOGIC;
    SIGNAL S4471 : STD_LOGIC;
    SIGNAL S4472 : STD_LOGIC;
    SIGNAL S4473 : STD_LOGIC;
    SIGNAL S4474 : STD_LOGIC;
    SIGNAL S4475 : STD_LOGIC;
    SIGNAL S4476 : STD_LOGIC;
    SIGNAL S4477 : STD_LOGIC;
    SIGNAL S4478 : STD_LOGIC;
    SIGNAL S4479 : STD_LOGIC;
    SIGNAL S4480 : STD_LOGIC;
    SIGNAL S4481 : STD_LOGIC;
    SIGNAL S4482 : STD_LOGIC;
    SIGNAL S4483 : STD_LOGIC;
    SIGNAL S4484 : STD_LOGIC;
    SIGNAL S4485 : STD_LOGIC;
    SIGNAL S4486 : STD_LOGIC;
    SIGNAL S4487 : STD_LOGIC;
    SIGNAL S4488 : STD_LOGIC;
    SIGNAL S4489 : STD_LOGIC;
    SIGNAL S4490 : STD_LOGIC;
    SIGNAL S4491 : STD_LOGIC;
    SIGNAL S4492 : STD_LOGIC;
    SIGNAL S4493 : STD_LOGIC;
    SIGNAL S4494 : STD_LOGIC;
    SIGNAL S4495 : STD_LOGIC;
    SIGNAL S4496 : STD_LOGIC;
    SIGNAL S4497 : STD_LOGIC;
    SIGNAL S4498 : STD_LOGIC;
    SIGNAL S4499 : STD_LOGIC;
    SIGNAL S4500 : STD_LOGIC;
    SIGNAL S4501 : STD_LOGIC;
    SIGNAL S4502 : STD_LOGIC;
    SIGNAL S4503 : STD_LOGIC;
    SIGNAL S4504 : STD_LOGIC;
    SIGNAL S4505 : STD_LOGIC;
    SIGNAL S4506 : STD_LOGIC;
    SIGNAL S4507 : STD_LOGIC;
    SIGNAL S4508 : STD_LOGIC;
    SIGNAL S4509 : STD_LOGIC;
    SIGNAL S4510 : STD_LOGIC;
    SIGNAL S4511 : STD_LOGIC;
    SIGNAL S4512 : STD_LOGIC;
    SIGNAL S4513 : STD_LOGIC;
    SIGNAL S4514 : STD_LOGIC;
    SIGNAL S4515 : STD_LOGIC;
    SIGNAL S4516 : STD_LOGIC;
    SIGNAL S4517 : STD_LOGIC;
    SIGNAL S4518 : STD_LOGIC;
    SIGNAL S4519 : STD_LOGIC;
    SIGNAL S4520 : STD_LOGIC;
    SIGNAL S4521 : STD_LOGIC;
    SIGNAL S4522 : STD_LOGIC;
    SIGNAL S4523 : STD_LOGIC;
    SIGNAL S4524 : STD_LOGIC;
    SIGNAL S4525 : STD_LOGIC;
    SIGNAL S4526 : STD_LOGIC;
    SIGNAL S4527 : STD_LOGIC;
    SIGNAL S4528 : STD_LOGIC;
    SIGNAL S4529 : STD_LOGIC;
    SIGNAL S4530 : STD_LOGIC;
    SIGNAL S4531 : STD_LOGIC;
    SIGNAL S4532 : STD_LOGIC;
    SIGNAL S4533 : STD_LOGIC;
    SIGNAL S4534 : STD_LOGIC;
    SIGNAL S4535 : STD_LOGIC;
    SIGNAL S4536 : STD_LOGIC;
    SIGNAL S4537 : STD_LOGIC;
    SIGNAL S4538 : STD_LOGIC;
    SIGNAL S4539 : STD_LOGIC;
    SIGNAL S4540 : STD_LOGIC;
    SIGNAL S4541 : STD_LOGIC;
    SIGNAL S4542 : STD_LOGIC;
    SIGNAL S4543 : STD_LOGIC;
    SIGNAL S4544 : STD_LOGIC;
    SIGNAL S4545 : STD_LOGIC;
    SIGNAL S4546 : STD_LOGIC;
    SIGNAL S4547 : STD_LOGIC;
    SIGNAL S4548 : STD_LOGIC;
    SIGNAL S4549 : STD_LOGIC;
    SIGNAL S4550 : STD_LOGIC;
    SIGNAL S4551 : STD_LOGIC;
    SIGNAL S4552 : STD_LOGIC;
    SIGNAL S4553 : STD_LOGIC;
    SIGNAL S4554 : STD_LOGIC;
    SIGNAL S4555 : STD_LOGIC;
    SIGNAL S4556 : STD_LOGIC;
    SIGNAL S4557 : STD_LOGIC;
    SIGNAL S4558 : STD_LOGIC;
    SIGNAL S4559 : STD_LOGIC;
    SIGNAL S4560 : STD_LOGIC;
    SIGNAL S4561 : STD_LOGIC;
    SIGNAL S4562 : STD_LOGIC;
    SIGNAL S4563 : STD_LOGIC;
    SIGNAL S4564 : STD_LOGIC;
    SIGNAL S4565 : STD_LOGIC;
    SIGNAL S4566 : STD_LOGIC;
    SIGNAL S4567 : STD_LOGIC;
    SIGNAL S4568 : STD_LOGIC;
    SIGNAL S4569 : STD_LOGIC;
    SIGNAL S4570 : STD_LOGIC;
    SIGNAL S4571 : STD_LOGIC;
    SIGNAL S4572 : STD_LOGIC;
    SIGNAL S4573 : STD_LOGIC;
    SIGNAL S4574 : STD_LOGIC;
    SIGNAL S4575 : STD_LOGIC;
    SIGNAL S4576 : STD_LOGIC;
    SIGNAL S4577 : STD_LOGIC;
    SIGNAL S4578 : STD_LOGIC;
    SIGNAL S4579 : STD_LOGIC;
    SIGNAL S4580 : STD_LOGIC;
    SIGNAL S4581 : STD_LOGIC;
    SIGNAL S4582 : STD_LOGIC;
    SIGNAL S4583 : STD_LOGIC;
    SIGNAL S4584 : STD_LOGIC;
    SIGNAL S4585 : STD_LOGIC;
    SIGNAL S4586 : STD_LOGIC;
    SIGNAL S4587 : STD_LOGIC;
    SIGNAL S4588 : STD_LOGIC;
    SIGNAL S4589 : STD_LOGIC;
    SIGNAL S4590 : STD_LOGIC;
    SIGNAL S4591 : STD_LOGIC;
    SIGNAL S4592 : STD_LOGIC;
    SIGNAL S4593 : STD_LOGIC;
    SIGNAL S4594 : STD_LOGIC;
    SIGNAL S4595 : STD_LOGIC;
    SIGNAL S4596 : STD_LOGIC;
    SIGNAL S4597 : STD_LOGIC;
    SIGNAL S4598 : STD_LOGIC;
    SIGNAL S4599 : STD_LOGIC;
    SIGNAL S4600 : STD_LOGIC;
    SIGNAL S4601 : STD_LOGIC;
    SIGNAL S4602 : STD_LOGIC;
    SIGNAL S4603 : STD_LOGIC;
    SIGNAL S4604 : STD_LOGIC;
    SIGNAL S4605 : STD_LOGIC;
    SIGNAL S4606 : STD_LOGIC;
    SIGNAL S4607 : STD_LOGIC;
    SIGNAL S4608 : STD_LOGIC;
    SIGNAL S4609 : STD_LOGIC;
    SIGNAL S4610 : STD_LOGIC;
    SIGNAL S4611 : STD_LOGIC;
    SIGNAL S4612 : STD_LOGIC;
    SIGNAL S4613 : STD_LOGIC;
    SIGNAL S4614 : STD_LOGIC;
    SIGNAL S4615 : STD_LOGIC;
    SIGNAL S4616 : STD_LOGIC;
    SIGNAL S4617 : STD_LOGIC;
    SIGNAL S4618 : STD_LOGIC;
    SIGNAL S4619 : STD_LOGIC;
    SIGNAL S4620 : STD_LOGIC;
    SIGNAL S4621 : STD_LOGIC;
    SIGNAL S4622 : STD_LOGIC;
    SIGNAL S4623 : STD_LOGIC;
    SIGNAL S4624 : STD_LOGIC;
    SIGNAL S4625 : STD_LOGIC;
    SIGNAL S4626 : STD_LOGIC;
    SIGNAL S4627 : STD_LOGIC;
    SIGNAL S4628 : STD_LOGIC;
    SIGNAL S4629 : STD_LOGIC;
    SIGNAL S4630 : STD_LOGIC;
    SIGNAL S4631 : STD_LOGIC;
    SIGNAL S4632 : STD_LOGIC;
    SIGNAL S4633 : STD_LOGIC;
    SIGNAL S4634 : STD_LOGIC;
    SIGNAL S4635 : STD_LOGIC;
    SIGNAL S4636 : STD_LOGIC;
    SIGNAL S4637 : STD_LOGIC;
    SIGNAL S4638 : STD_LOGIC;
    SIGNAL S4639 : STD_LOGIC;
    SIGNAL S4640 : STD_LOGIC;
    SIGNAL S4641 : STD_LOGIC;
    SIGNAL S4642 : STD_LOGIC;
    SIGNAL S4643 : STD_LOGIC;
    SIGNAL S4644 : STD_LOGIC;
    SIGNAL S4645 : STD_LOGIC;
    SIGNAL S4646 : STD_LOGIC;
    SIGNAL S4647 : STD_LOGIC;
    SIGNAL S4648 : STD_LOGIC;
    SIGNAL S4649 : STD_LOGIC;
    SIGNAL S4650 : STD_LOGIC;
    SIGNAL S4651 : STD_LOGIC;
    SIGNAL S4652 : STD_LOGIC;
    SIGNAL S4653 : STD_LOGIC;
    SIGNAL S4654 : STD_LOGIC;
    SIGNAL S4655 : STD_LOGIC;
    SIGNAL S4656 : STD_LOGIC;
    SIGNAL S4657 : STD_LOGIC;
    SIGNAL S4658 : STD_LOGIC;
    SIGNAL S4659 : STD_LOGIC;
    SIGNAL S4660 : STD_LOGIC;
    SIGNAL S4661 : STD_LOGIC;
    SIGNAL S4662 : STD_LOGIC;
    SIGNAL S4663 : STD_LOGIC;
    SIGNAL S4664 : STD_LOGIC;
    SIGNAL S4665 : STD_LOGIC;
    SIGNAL S4666 : STD_LOGIC;
    SIGNAL S4667 : STD_LOGIC;
    SIGNAL S4668 : STD_LOGIC;
    SIGNAL S4669 : STD_LOGIC;
    SIGNAL S4670 : STD_LOGIC;
    SIGNAL S4671 : STD_LOGIC;
    SIGNAL S4672 : STD_LOGIC;
    SIGNAL S4673 : STD_LOGIC;
    SIGNAL S4674 : STD_LOGIC;
    SIGNAL S4675 : STD_LOGIC;
    SIGNAL S4676 : STD_LOGIC;
    SIGNAL S4677 : STD_LOGIC;
    SIGNAL S4678 : STD_LOGIC;
    SIGNAL S4679 : STD_LOGIC;
    SIGNAL S4680 : STD_LOGIC;
    SIGNAL S4681 : STD_LOGIC;
    SIGNAL S4682 : STD_LOGIC;
    SIGNAL S4683 : STD_LOGIC;
    SIGNAL S4684 : STD_LOGIC;
    SIGNAL S4685 : STD_LOGIC;
    SIGNAL S4686 : STD_LOGIC;
    SIGNAL S4687 : STD_LOGIC;
    SIGNAL S4688 : STD_LOGIC;
    SIGNAL S4689 : STD_LOGIC;
    SIGNAL S4690 : STD_LOGIC;
    SIGNAL S4691 : STD_LOGIC;
    SIGNAL S4692 : STD_LOGIC;
    SIGNAL S4693 : STD_LOGIC;
    SIGNAL S4694 : STD_LOGIC;
    SIGNAL S4695 : STD_LOGIC;
    SIGNAL S4696 : STD_LOGIC;
    SIGNAL S4697 : STD_LOGIC;
    SIGNAL S4698 : STD_LOGIC;
    SIGNAL S4699 : STD_LOGIC;
    SIGNAL S4700 : STD_LOGIC;
    SIGNAL S4701 : STD_LOGIC;
    SIGNAL S4702 : STD_LOGIC;
    SIGNAL S4703 : STD_LOGIC;
    SIGNAL S4704 : STD_LOGIC;
    SIGNAL S4705 : STD_LOGIC;
    SIGNAL S4706 : STD_LOGIC;
    SIGNAL S4707 : STD_LOGIC;
    SIGNAL S4708 : STD_LOGIC;
    SIGNAL S4709 : STD_LOGIC;
    SIGNAL S4710 : STD_LOGIC;
    SIGNAL S4711 : STD_LOGIC;
    SIGNAL S4712 : STD_LOGIC;
    SIGNAL S4713 : STD_LOGIC;
    SIGNAL S4714 : STD_LOGIC;
    SIGNAL S4715 : STD_LOGIC;
    SIGNAL S4716 : STD_LOGIC;
    SIGNAL S4717 : STD_LOGIC;
    SIGNAL S4718 : STD_LOGIC;
    SIGNAL S4719 : STD_LOGIC;
    SIGNAL S4720 : STD_LOGIC;
    SIGNAL S4721 : STD_LOGIC;
    SIGNAL S4722 : STD_LOGIC;
    SIGNAL S4723 : STD_LOGIC;
    SIGNAL S4724 : STD_LOGIC;
    SIGNAL S4725 : STD_LOGIC;
    SIGNAL S4726 : STD_LOGIC;
    SIGNAL S4727 : STD_LOGIC;
    SIGNAL S4728 : STD_LOGIC;
    SIGNAL S4729 : STD_LOGIC;
    SIGNAL S4730 : STD_LOGIC;
    SIGNAL S4731 : STD_LOGIC;
    SIGNAL S4732 : STD_LOGIC;
    SIGNAL S4733 : STD_LOGIC;
    SIGNAL S4734 : STD_LOGIC;
    SIGNAL S4735 : STD_LOGIC;
    SIGNAL S4736 : STD_LOGIC;
    SIGNAL S4737 : STD_LOGIC;
    SIGNAL S4738 : STD_LOGIC;
    SIGNAL S4739 : STD_LOGIC;
    SIGNAL S4740 : STD_LOGIC;
    SIGNAL S4741 : STD_LOGIC;
    SIGNAL S4742 : STD_LOGIC;
    SIGNAL S4743 : STD_LOGIC;
    SIGNAL S4744 : STD_LOGIC;
    SIGNAL S4745 : STD_LOGIC;
    SIGNAL S4746 : STD_LOGIC;
    SIGNAL S4747 : STD_LOGIC;
    SIGNAL S4748 : STD_LOGIC;
    SIGNAL S4749 : STD_LOGIC;
    SIGNAL S4750 : STD_LOGIC;
    SIGNAL S4751 : STD_LOGIC;
    SIGNAL S4752 : STD_LOGIC;
    SIGNAL S4753 : STD_LOGIC;
    SIGNAL S4754 : STD_LOGIC;
    SIGNAL S4755 : STD_LOGIC;
    SIGNAL S4756 : STD_LOGIC;
    SIGNAL S4757 : STD_LOGIC;
    SIGNAL S4758 : STD_LOGIC;
    SIGNAL S4759 : STD_LOGIC;
    SIGNAL S4760 : STD_LOGIC;
    SIGNAL S4761 : STD_LOGIC;
    SIGNAL S4762 : STD_LOGIC;
    SIGNAL S4763 : STD_LOGIC;
    SIGNAL S4764 : STD_LOGIC;
    SIGNAL S4765 : STD_LOGIC;
    SIGNAL S4766 : STD_LOGIC;
    SIGNAL S4767 : STD_LOGIC;
    SIGNAL S4768 : STD_LOGIC;
    SIGNAL S4769 : STD_LOGIC;
    SIGNAL S4770 : STD_LOGIC;
    SIGNAL S4771 : STD_LOGIC;
    SIGNAL S4772 : STD_LOGIC;
    SIGNAL S4773 : STD_LOGIC;
    SIGNAL S4774 : STD_LOGIC;
    SIGNAL S4775 : STD_LOGIC;
    SIGNAL S4776 : STD_LOGIC;
    SIGNAL S4777 : STD_LOGIC;
    SIGNAL S4778 : STD_LOGIC;
    SIGNAL S4779 : STD_LOGIC;
    SIGNAL S4780 : STD_LOGIC;
    SIGNAL S4781 : STD_LOGIC;
    SIGNAL S4782 : STD_LOGIC;
    SIGNAL S4783 : STD_LOGIC;
    SIGNAL S4784 : STD_LOGIC;
    SIGNAL S4785 : STD_LOGIC;
    SIGNAL S4786 : STD_LOGIC;
    SIGNAL S4787 : STD_LOGIC;
    SIGNAL S4788 : STD_LOGIC;
    SIGNAL S4789 : STD_LOGIC;
    SIGNAL S4790 : STD_LOGIC;
    SIGNAL S4791 : STD_LOGIC;
    SIGNAL S4792 : STD_LOGIC;
    SIGNAL S4793 : STD_LOGIC;
    SIGNAL S4794 : STD_LOGIC;
    SIGNAL S4795 : STD_LOGIC;
    SIGNAL S4796 : STD_LOGIC;
    SIGNAL S4797 : STD_LOGIC;
    SIGNAL S4798 : STD_LOGIC;
    SIGNAL S4799 : STD_LOGIC;
    SIGNAL S4800 : STD_LOGIC;
    SIGNAL S4801 : STD_LOGIC;
    SIGNAL S4802 : STD_LOGIC;
    SIGNAL S4803 : STD_LOGIC;
    SIGNAL S4804 : STD_LOGIC;
    SIGNAL S4805 : STD_LOGIC;
    SIGNAL S4806 : STD_LOGIC;
    SIGNAL S4807 : STD_LOGIC;
    SIGNAL S4808 : STD_LOGIC;
    SIGNAL S4809 : STD_LOGIC;
    SIGNAL S4810 : STD_LOGIC;
    SIGNAL S4811 : STD_LOGIC;
    SIGNAL S4812 : STD_LOGIC;
    SIGNAL S4813 : STD_LOGIC;
    SIGNAL S4814 : STD_LOGIC;
    SIGNAL S4815 : STD_LOGIC;
    SIGNAL S4816 : STD_LOGIC;
    SIGNAL S4817 : STD_LOGIC;
    SIGNAL S4818 : STD_LOGIC;
    SIGNAL S4819 : STD_LOGIC;
    SIGNAL S4820 : STD_LOGIC;
    SIGNAL S4821 : STD_LOGIC;
    SIGNAL S4822 : STD_LOGIC;
    SIGNAL S4823 : STD_LOGIC;
    SIGNAL S4824 : STD_LOGIC;
    SIGNAL S4825 : STD_LOGIC;
    SIGNAL S4826 : STD_LOGIC;
    SIGNAL S4827 : STD_LOGIC;
    SIGNAL S4828 : STD_LOGIC;
    SIGNAL S4829 : STD_LOGIC;
    SIGNAL S4830 : STD_LOGIC;
    SIGNAL S4831 : STD_LOGIC;
    SIGNAL S4832 : STD_LOGIC;
    SIGNAL S4833 : STD_LOGIC;
    SIGNAL S4834 : STD_LOGIC;
    SIGNAL S4835 : STD_LOGIC;
    SIGNAL S4836 : STD_LOGIC;
    SIGNAL S4837 : STD_LOGIC;
    SIGNAL S4838 : STD_LOGIC;
    SIGNAL S4839 : STD_LOGIC;
    SIGNAL S4840 : STD_LOGIC;
    SIGNAL S4841 : STD_LOGIC;
    SIGNAL S4842 : STD_LOGIC;
    SIGNAL S4843 : STD_LOGIC;
    SIGNAL S4844 : STD_LOGIC;
    SIGNAL S4845 : STD_LOGIC;
    SIGNAL S4846 : STD_LOGIC;
    SIGNAL S4847 : STD_LOGIC;
    SIGNAL S4848 : STD_LOGIC;
    SIGNAL S4849 : STD_LOGIC;
    SIGNAL S4850 : STD_LOGIC;
    SIGNAL S4851 : STD_LOGIC;
    SIGNAL S4852 : STD_LOGIC;
    SIGNAL S4853 : STD_LOGIC;
    SIGNAL S4854 : STD_LOGIC;
    SIGNAL S4855 : STD_LOGIC;
    SIGNAL S4856 : STD_LOGIC;
    SIGNAL S4857 : STD_LOGIC;
    SIGNAL S4858 : STD_LOGIC;
    SIGNAL S4859 : STD_LOGIC;
    SIGNAL S4860 : STD_LOGIC;
    SIGNAL S4861 : STD_LOGIC;
    SIGNAL S4862 : STD_LOGIC;
    SIGNAL S4863 : STD_LOGIC;
    SIGNAL S4864 : STD_LOGIC;
    SIGNAL S4865 : STD_LOGIC;
    SIGNAL S4866 : STD_LOGIC;
    SIGNAL S4867 : STD_LOGIC;
    SIGNAL S4868 : STD_LOGIC;
    SIGNAL S4869 : STD_LOGIC;
    SIGNAL S4870 : STD_LOGIC;
    SIGNAL S4871 : STD_LOGIC;
    SIGNAL S4872 : STD_LOGIC;
    SIGNAL S4873 : STD_LOGIC;
    SIGNAL S4874 : STD_LOGIC;
    SIGNAL S4875 : STD_LOGIC;
    SIGNAL S4876 : STD_LOGIC;
    SIGNAL S4877 : STD_LOGIC;
    SIGNAL S4878 : STD_LOGIC;
    SIGNAL S4879 : STD_LOGIC;
    SIGNAL S4880 : STD_LOGIC;
    SIGNAL S4881 : STD_LOGIC;
    SIGNAL S4882 : STD_LOGIC;
    SIGNAL S4883 : STD_LOGIC;
    SIGNAL S4884 : STD_LOGIC;
    SIGNAL S4885 : STD_LOGIC;
    SIGNAL S4886 : STD_LOGIC;
    SIGNAL S4887 : STD_LOGIC;
    SIGNAL S4888 : STD_LOGIC;
    SIGNAL S4889 : STD_LOGIC;
    SIGNAL S4890 : STD_LOGIC;
    SIGNAL S4891 : STD_LOGIC;
    SIGNAL S4892 : STD_LOGIC;
    SIGNAL S4893 : STD_LOGIC;
    SIGNAL S4894 : STD_LOGIC;
    SIGNAL S4895 : STD_LOGIC;
    SIGNAL S4896 : STD_LOGIC;
    SIGNAL S4897 : STD_LOGIC;
    SIGNAL S4898 : STD_LOGIC;
    SIGNAL S4899 : STD_LOGIC;
    SIGNAL S4900 : STD_LOGIC;
    SIGNAL S4901 : STD_LOGIC;
    SIGNAL S4902 : STD_LOGIC;
    SIGNAL S4903 : STD_LOGIC;
    SIGNAL S4904 : STD_LOGIC;
    SIGNAL S4905 : STD_LOGIC;
    SIGNAL S4906 : STD_LOGIC;
    SIGNAL S4907 : STD_LOGIC;
    SIGNAL S4908 : STD_LOGIC;
    SIGNAL S4909 : STD_LOGIC;
    SIGNAL S4910 : STD_LOGIC;
    SIGNAL S4911 : STD_LOGIC;
    SIGNAL S4912 : STD_LOGIC;
    SIGNAL S4913 : STD_LOGIC;
    SIGNAL S4914 : STD_LOGIC;
    SIGNAL S4915 : STD_LOGIC;
    SIGNAL S4916 : STD_LOGIC;
    SIGNAL S4917 : STD_LOGIC;
    SIGNAL S4918 : STD_LOGIC;
    SIGNAL S4919 : STD_LOGIC;
    SIGNAL S4920 : STD_LOGIC;
    SIGNAL S4921 : STD_LOGIC;
    SIGNAL S4922 : STD_LOGIC;
    SIGNAL S4923 : STD_LOGIC;
    SIGNAL S4924 : STD_LOGIC;
    SIGNAL S4925 : STD_LOGIC;
    SIGNAL S4926 : STD_LOGIC;
    SIGNAL S4927 : STD_LOGIC;
    SIGNAL S4928 : STD_LOGIC;
    SIGNAL S4929 : STD_LOGIC;
    SIGNAL S4930 : STD_LOGIC;
    SIGNAL S4931 : STD_LOGIC;
    SIGNAL S4932 : STD_LOGIC;
    SIGNAL S4933 : STD_LOGIC;
    SIGNAL S4934 : STD_LOGIC;
    SIGNAL S4935 : STD_LOGIC;
    SIGNAL S4936 : STD_LOGIC;
    SIGNAL S4937 : STD_LOGIC;
    SIGNAL S4938 : STD_LOGIC;
    SIGNAL S4939 : STD_LOGIC;
    SIGNAL S4940 : STD_LOGIC;
    SIGNAL S4941 : STD_LOGIC;
    SIGNAL S4942 : STD_LOGIC;
    SIGNAL S4943 : STD_LOGIC;
    SIGNAL S4944 : STD_LOGIC;
    SIGNAL S4945 : STD_LOGIC;
    SIGNAL S4946 : STD_LOGIC;
    SIGNAL S4947 : STD_LOGIC;
    SIGNAL S4948 : STD_LOGIC;
    SIGNAL S4949 : STD_LOGIC;
    SIGNAL S4950 : STD_LOGIC;
    SIGNAL S4951 : STD_LOGIC;
    SIGNAL S4952 : STD_LOGIC;
    SIGNAL S4953 : STD_LOGIC;
    SIGNAL S4954 : STD_LOGIC;
    SIGNAL S4955 : STD_LOGIC;
    SIGNAL S4956 : STD_LOGIC;
    SIGNAL S4957 : STD_LOGIC;
    SIGNAL S4958 : STD_LOGIC;
    SIGNAL S4959 : STD_LOGIC;
    SIGNAL S4960 : STD_LOGIC;
    SIGNAL S4961 : STD_LOGIC;
    SIGNAL S4962 : STD_LOGIC;
    SIGNAL S4963 : STD_LOGIC;
    SIGNAL S4964 : STD_LOGIC;
    SIGNAL S4965 : STD_LOGIC;
    SIGNAL S4966 : STD_LOGIC;
    SIGNAL S4967 : STD_LOGIC;
    SIGNAL S4968 : STD_LOGIC;
    SIGNAL S4969 : STD_LOGIC;
    SIGNAL S4970 : STD_LOGIC;
    SIGNAL S4971 : STD_LOGIC;
    SIGNAL S4972 : STD_LOGIC;
    SIGNAL S4973 : STD_LOGIC;
    SIGNAL S4974 : STD_LOGIC;
    SIGNAL S4975 : STD_LOGIC;
    SIGNAL S4976 : STD_LOGIC;
    SIGNAL S4977 : STD_LOGIC;
    SIGNAL S4978 : STD_LOGIC;
    SIGNAL S4979 : STD_LOGIC;
    SIGNAL S4980 : STD_LOGIC;
    SIGNAL S4981 : STD_LOGIC;
    SIGNAL S4982 : STD_LOGIC;
    SIGNAL S4983 : STD_LOGIC;
    SIGNAL S4984 : STD_LOGIC;
    SIGNAL S4985 : STD_LOGIC;
    SIGNAL S4986 : STD_LOGIC;
    SIGNAL S4987 : STD_LOGIC;
    SIGNAL S4988 : STD_LOGIC;
    SIGNAL S4989 : STD_LOGIC;
    SIGNAL S4990 : STD_LOGIC;
    SIGNAL S4991 : STD_LOGIC;
    SIGNAL S4992 : STD_LOGIC;
    SIGNAL S4993 : STD_LOGIC;
    SIGNAL S4994 : STD_LOGIC;
    SIGNAL S4995 : STD_LOGIC;
    SIGNAL S4996 : STD_LOGIC;
    SIGNAL S4997 : STD_LOGIC;
    SIGNAL S4998 : STD_LOGIC;
    SIGNAL S4999 : STD_LOGIC;
    SIGNAL S5000 : STD_LOGIC;
    SIGNAL S5001 : STD_LOGIC;
    SIGNAL S5002 : STD_LOGIC;
    SIGNAL S5003 : STD_LOGIC;
    SIGNAL S5004 : STD_LOGIC;
    SIGNAL S5005 : STD_LOGIC;
    SIGNAL S5006 : STD_LOGIC;
    SIGNAL S5007 : STD_LOGIC;
    SIGNAL S5008 : STD_LOGIC;
    SIGNAL S5009 : STD_LOGIC;
    SIGNAL S5010 : STD_LOGIC;
    SIGNAL S5011 : STD_LOGIC;
    SIGNAL S5012 : STD_LOGIC;
    SIGNAL S5013 : STD_LOGIC;
    SIGNAL S5014 : STD_LOGIC;
    SIGNAL S5015 : STD_LOGIC;
    SIGNAL S5016 : STD_LOGIC;
    SIGNAL S5017 : STD_LOGIC;
    SIGNAL S5018 : STD_LOGIC;
    SIGNAL S5019 : STD_LOGIC;
    SIGNAL S5020 : STD_LOGIC;
    SIGNAL S5021 : STD_LOGIC;
    SIGNAL S5022 : STD_LOGIC;
    SIGNAL S5023 : STD_LOGIC;
    SIGNAL S5024 : STD_LOGIC;
    SIGNAL S5025 : STD_LOGIC;
    SIGNAL S5026 : STD_LOGIC;
    SIGNAL S5027 : STD_LOGIC;
    SIGNAL S5028 : STD_LOGIC;
    SIGNAL S5029 : STD_LOGIC;
    SIGNAL S5030 : STD_LOGIC;
    SIGNAL S5031 : STD_LOGIC;
    SIGNAL S5032 : STD_LOGIC;
    SIGNAL S5033 : STD_LOGIC;
    SIGNAL S5034 : STD_LOGIC;
    SIGNAL S5035 : STD_LOGIC;
    SIGNAL S5036 : STD_LOGIC;
    SIGNAL S5037 : STD_LOGIC;
    SIGNAL S5038 : STD_LOGIC;
    SIGNAL S5039 : STD_LOGIC;
    SIGNAL S5040 : STD_LOGIC;
    SIGNAL S5041 : STD_LOGIC;
    SIGNAL S5042 : STD_LOGIC;
    SIGNAL S5043 : STD_LOGIC;
    SIGNAL S5044 : STD_LOGIC;
    SIGNAL S5045 : STD_LOGIC;
    SIGNAL S5046 : STD_LOGIC;
    SIGNAL S5047 : STD_LOGIC;
    SIGNAL S5048 : STD_LOGIC;
    SIGNAL S5049 : STD_LOGIC;
    SIGNAL S5050 : STD_LOGIC;
    SIGNAL S5051 : STD_LOGIC;
    SIGNAL S5052 : STD_LOGIC;
    SIGNAL S5053 : STD_LOGIC;
    SIGNAL S5054 : STD_LOGIC;
    SIGNAL S5055 : STD_LOGIC;
    SIGNAL S5056 : STD_LOGIC;
    SIGNAL S5057 : STD_LOGIC;
    SIGNAL S5058 : STD_LOGIC;
    SIGNAL S5059 : STD_LOGIC;
    SIGNAL S5060 : STD_LOGIC;
    SIGNAL S5061 : STD_LOGIC;
    SIGNAL S5062 : STD_LOGIC;
    SIGNAL S5063 : STD_LOGIC;
    SIGNAL S5064 : STD_LOGIC;
    SIGNAL S5065 : STD_LOGIC;
    SIGNAL S5066 : STD_LOGIC;
    SIGNAL S5067 : STD_LOGIC;
    SIGNAL S5068 : STD_LOGIC;
    SIGNAL S5069 : STD_LOGIC;
    SIGNAL S5070 : STD_LOGIC;
    SIGNAL S5071 : STD_LOGIC;
    SIGNAL S5072 : STD_LOGIC;
    SIGNAL S5073 : STD_LOGIC;
    SIGNAL S5074 : STD_LOGIC;
    SIGNAL S5075 : STD_LOGIC;
    SIGNAL S5076 : STD_LOGIC;
    SIGNAL S5077 : STD_LOGIC;
    SIGNAL S5078 : STD_LOGIC;
    SIGNAL S5079 : STD_LOGIC;
    SIGNAL S5080 : STD_LOGIC;
    SIGNAL S5081 : STD_LOGIC;
    SIGNAL S5082 : STD_LOGIC;
    SIGNAL S5083 : STD_LOGIC;
    SIGNAL S5084 : STD_LOGIC;
    SIGNAL S5085 : STD_LOGIC;
    SIGNAL S5086 : STD_LOGIC;
    SIGNAL S5087 : STD_LOGIC;
    SIGNAL S5088 : STD_LOGIC;
    SIGNAL S5089 : STD_LOGIC;
    SIGNAL S5090 : STD_LOGIC;
    SIGNAL S5091 : STD_LOGIC;
    SIGNAL S5092 : STD_LOGIC;
    SIGNAL S5093 : STD_LOGIC;
    SIGNAL S5094 : STD_LOGIC;
    SIGNAL S5095 : STD_LOGIC;
    SIGNAL S5096 : STD_LOGIC;
    SIGNAL S5097 : STD_LOGIC;
    SIGNAL S5098 : STD_LOGIC;
    SIGNAL S5099 : STD_LOGIC;
    SIGNAL S5100 : STD_LOGIC;
    SIGNAL S5101 : STD_LOGIC;
    SIGNAL S5102 : STD_LOGIC;
    SIGNAL S5103 : STD_LOGIC;
    SIGNAL S5104 : STD_LOGIC;
    SIGNAL S5105 : STD_LOGIC;
    SIGNAL S5106 : STD_LOGIC;
    SIGNAL S5107 : STD_LOGIC;
    SIGNAL S5108 : STD_LOGIC;
    SIGNAL S5109 : STD_LOGIC;
    SIGNAL S5110 : STD_LOGIC;
    SIGNAL S5111 : STD_LOGIC;
    SIGNAL S5112 : STD_LOGIC;
    SIGNAL S5113 : STD_LOGIC;
    SIGNAL S5114 : STD_LOGIC;
    SIGNAL S5115 : STD_LOGIC;
    SIGNAL S5116 : STD_LOGIC;
    SIGNAL S5117 : STD_LOGIC;
    SIGNAL S5118 : STD_LOGIC;
    SIGNAL S5119 : STD_LOGIC;
    SIGNAL S5120 : STD_LOGIC;
    SIGNAL S5121 : STD_LOGIC;
    SIGNAL S5122 : STD_LOGIC;
    SIGNAL S5123 : STD_LOGIC;
    SIGNAL S5124 : STD_LOGIC;
    SIGNAL S5125 : STD_LOGIC;
    SIGNAL S5126 : STD_LOGIC;
    SIGNAL S5127 : STD_LOGIC;
    SIGNAL S5128 : STD_LOGIC;
    SIGNAL S5129 : STD_LOGIC;
    SIGNAL S5130 : STD_LOGIC;
    SIGNAL S5131 : STD_LOGIC;
    SIGNAL S5132 : STD_LOGIC;
    SIGNAL S5133 : STD_LOGIC;
    SIGNAL S5134 : STD_LOGIC;
    SIGNAL S5135 : STD_LOGIC;
    SIGNAL S5136 : STD_LOGIC;
    SIGNAL S5137 : STD_LOGIC;
    SIGNAL S5138 : STD_LOGIC;
    SIGNAL S5139 : STD_LOGIC;
    SIGNAL S5140 : STD_LOGIC;
    SIGNAL S5141 : STD_LOGIC;
    SIGNAL S5142 : STD_LOGIC;
    SIGNAL S5143 : STD_LOGIC;
    SIGNAL S5144 : STD_LOGIC;
    SIGNAL S5145 : STD_LOGIC;
    SIGNAL S5146 : STD_LOGIC;
    SIGNAL S5147 : STD_LOGIC;
    SIGNAL S5148 : STD_LOGIC;
    SIGNAL S5149 : STD_LOGIC;
    SIGNAL S5150 : STD_LOGIC;
    SIGNAL S5151 : STD_LOGIC;
    SIGNAL S5152 : STD_LOGIC;
    SIGNAL S5153 : STD_LOGIC;
    SIGNAL S5154 : STD_LOGIC;
    SIGNAL S5155 : STD_LOGIC;
    SIGNAL S5156 : STD_LOGIC;
    SIGNAL S5157 : STD_LOGIC;
    SIGNAL S5158 : STD_LOGIC;
    SIGNAL S5159 : STD_LOGIC;
    SIGNAL S5160 : STD_LOGIC;
    SIGNAL S5161 : STD_LOGIC;
    SIGNAL S5162 : STD_LOGIC;
    SIGNAL S5163 : STD_LOGIC;
    SIGNAL S5164 : STD_LOGIC;
    SIGNAL S5165 : STD_LOGIC;
    SIGNAL S5166 : STD_LOGIC;
    SIGNAL S5167 : STD_LOGIC;
    SIGNAL S5168 : STD_LOGIC;
    SIGNAL S5169 : STD_LOGIC;
    SIGNAL S5170 : STD_LOGIC;
    SIGNAL S5171 : STD_LOGIC;
    SIGNAL S5172 : STD_LOGIC;
    SIGNAL S5173 : STD_LOGIC;
    SIGNAL S5174 : STD_LOGIC;
    SIGNAL S5175 : STD_LOGIC;
    SIGNAL S5176 : STD_LOGIC;
    SIGNAL S5177 : STD_LOGIC;
    SIGNAL S5178 : STD_LOGIC;
    SIGNAL S5179 : STD_LOGIC;
    SIGNAL S5180 : STD_LOGIC;
    SIGNAL S5181 : STD_LOGIC;
    SIGNAL S5182 : STD_LOGIC;
    SIGNAL S5183 : STD_LOGIC;
    SIGNAL S5184 : STD_LOGIC;
    SIGNAL S5185 : STD_LOGIC;
    SIGNAL S5186 : STD_LOGIC;
    SIGNAL S5187 : STD_LOGIC;
    SIGNAL S5188 : STD_LOGIC;
    SIGNAL S5189 : STD_LOGIC;
    SIGNAL S5190 : STD_LOGIC;
    SIGNAL S5191 : STD_LOGIC;
    SIGNAL S5192 : STD_LOGIC;
    SIGNAL S5193 : STD_LOGIC;
    SIGNAL S5194 : STD_LOGIC;
    SIGNAL S5195 : STD_LOGIC;
    SIGNAL S5196 : STD_LOGIC;
    SIGNAL S5197 : STD_LOGIC;
    SIGNAL S5198 : STD_LOGIC;
    SIGNAL S5199 : STD_LOGIC;
    SIGNAL S5200 : STD_LOGIC;
    SIGNAL S5201 : STD_LOGIC;
    SIGNAL S5202 : STD_LOGIC;
    SIGNAL S5203 : STD_LOGIC;
    SIGNAL S5204 : STD_LOGIC;
    SIGNAL S5205 : STD_LOGIC;
    SIGNAL S5206 : STD_LOGIC;
    SIGNAL S5207 : STD_LOGIC;
    SIGNAL S5208 : STD_LOGIC;
    SIGNAL S5209 : STD_LOGIC;
    SIGNAL S5210 : STD_LOGIC;
    SIGNAL S5211 : STD_LOGIC;
    SIGNAL S5212 : STD_LOGIC;
    SIGNAL S5213 : STD_LOGIC;
    SIGNAL S5214 : STD_LOGIC;
    SIGNAL S5215 : STD_LOGIC;
    SIGNAL S5216 : STD_LOGIC;
    SIGNAL S5217 : STD_LOGIC;
    SIGNAL S5218 : STD_LOGIC;
    SIGNAL S5219 : STD_LOGIC;
    SIGNAL S5220 : STD_LOGIC;
    SIGNAL S5221 : STD_LOGIC;
    SIGNAL S5222 : STD_LOGIC;
    SIGNAL S5223 : STD_LOGIC;
    SIGNAL S5224 : STD_LOGIC;
    SIGNAL S5225 : STD_LOGIC;
    SIGNAL S5226 : STD_LOGIC;
    SIGNAL S5227 : STD_LOGIC;
    SIGNAL S5228 : STD_LOGIC;
    SIGNAL S5229 : STD_LOGIC;
    SIGNAL S5230 : STD_LOGIC;
    SIGNAL S5231 : STD_LOGIC;
    SIGNAL S5232 : STD_LOGIC;
    SIGNAL S5233 : STD_LOGIC;
    SIGNAL S5234 : STD_LOGIC;
    SIGNAL S5235 : STD_LOGIC;
    SIGNAL S5236 : STD_LOGIC;
    SIGNAL S5237 : STD_LOGIC;
    SIGNAL S5238 : STD_LOGIC;
    SIGNAL S5239 : STD_LOGIC;
    SIGNAL S5240 : STD_LOGIC;
    SIGNAL S5241 : STD_LOGIC;
    SIGNAL S5242 : STD_LOGIC;
    SIGNAL S5243 : STD_LOGIC;
    SIGNAL S5244 : STD_LOGIC;
    SIGNAL S5245 : STD_LOGIC;
    SIGNAL S5246 : STD_LOGIC;
    SIGNAL S5247 : STD_LOGIC;
    SIGNAL S5248 : STD_LOGIC;
    SIGNAL S5249 : STD_LOGIC;
    SIGNAL S5250 : STD_LOGIC;
    SIGNAL S5251 : STD_LOGIC;
    SIGNAL S5252 : STD_LOGIC;
    SIGNAL S5253 : STD_LOGIC;
    SIGNAL S5254 : STD_LOGIC;
    SIGNAL S5255 : STD_LOGIC;
    SIGNAL S5256 : STD_LOGIC;
    SIGNAL S5257 : STD_LOGIC;
    SIGNAL S5258 : STD_LOGIC;
    SIGNAL S5259 : STD_LOGIC;
    SIGNAL S5260 : STD_LOGIC;
    SIGNAL S5261 : STD_LOGIC;
    SIGNAL S5262 : STD_LOGIC;
    SIGNAL S5263 : STD_LOGIC;
    SIGNAL S5264 : STD_LOGIC;
    SIGNAL S5265 : STD_LOGIC;
    SIGNAL S5266 : STD_LOGIC;
    SIGNAL S5267 : STD_LOGIC;
    SIGNAL S5268 : STD_LOGIC;
    SIGNAL S5269 : STD_LOGIC;
    SIGNAL S5270 : STD_LOGIC;
    SIGNAL S5271 : STD_LOGIC;
    SIGNAL S5272 : STD_LOGIC;
    SIGNAL S5273 : STD_LOGIC;
    SIGNAL S5274 : STD_LOGIC;
    SIGNAL S5275 : STD_LOGIC;
    SIGNAL S5276 : STD_LOGIC;
    SIGNAL S5277 : STD_LOGIC;
    SIGNAL S5278 : STD_LOGIC;
    SIGNAL S5279 : STD_LOGIC;
    SIGNAL S5280 : STD_LOGIC;
    SIGNAL S5281 : STD_LOGIC;
    SIGNAL S5282 : STD_LOGIC;
    SIGNAL S5283 : STD_LOGIC;
    SIGNAL S5284 : STD_LOGIC;
    SIGNAL S5285 : STD_LOGIC;
    SIGNAL S5286 : STD_LOGIC;
    SIGNAL S5287 : STD_LOGIC;
    SIGNAL S5288 : STD_LOGIC;
    SIGNAL S5289 : STD_LOGIC;
    SIGNAL S5290 : STD_LOGIC;
    SIGNAL S5291 : STD_LOGIC;
    SIGNAL S5292 : STD_LOGIC;
    SIGNAL S5293 : STD_LOGIC;
    SIGNAL S5294 : STD_LOGIC;
    SIGNAL S5295 : STD_LOGIC;
    SIGNAL S5296 : STD_LOGIC;
    SIGNAL S5297 : STD_LOGIC;
    SIGNAL S5298 : STD_LOGIC;
    SIGNAL S5299 : STD_LOGIC;
    SIGNAL S5300 : STD_LOGIC;
    SIGNAL S5301 : STD_LOGIC;
    SIGNAL S5302 : STD_LOGIC;
    SIGNAL S5303 : STD_LOGIC;
    SIGNAL S5304 : STD_LOGIC;
    SIGNAL S5305 : STD_LOGIC;
    SIGNAL S5306 : STD_LOGIC;
    SIGNAL S5307 : STD_LOGIC;
    SIGNAL S5308 : STD_LOGIC;
    SIGNAL S5309 : STD_LOGIC;
    SIGNAL S5310 : STD_LOGIC;
    SIGNAL S5311 : STD_LOGIC;
    SIGNAL S5312 : STD_LOGIC;
    SIGNAL S5313 : STD_LOGIC;
    SIGNAL S5314 : STD_LOGIC;
    SIGNAL S5315 : STD_LOGIC;
    SIGNAL S5316 : STD_LOGIC;
    SIGNAL S5317 : STD_LOGIC;
    SIGNAL S5318 : STD_LOGIC;
    SIGNAL S5319 : STD_LOGIC;
    SIGNAL S5320 : STD_LOGIC;
    SIGNAL S5321 : STD_LOGIC;
    SIGNAL S5322 : STD_LOGIC;
    SIGNAL S5323 : STD_LOGIC;
    SIGNAL S5324 : STD_LOGIC;
    SIGNAL S5325 : STD_LOGIC;
    SIGNAL S5326 : STD_LOGIC;
    SIGNAL S5327 : STD_LOGIC;
    SIGNAL S5328 : STD_LOGIC;
    SIGNAL S5329 : STD_LOGIC;
    SIGNAL S5330 : STD_LOGIC;
    SIGNAL S5331 : STD_LOGIC;
    SIGNAL S5332 : STD_LOGIC;
    SIGNAL S5333 : STD_LOGIC;
    SIGNAL S5334 : STD_LOGIC;
    SIGNAL S5335 : STD_LOGIC;
    SIGNAL S5336 : STD_LOGIC;
    SIGNAL S5337 : STD_LOGIC;
    SIGNAL S5338 : STD_LOGIC;
    SIGNAL S5339 : STD_LOGIC;
    SIGNAL S5340 : STD_LOGIC;
    SIGNAL S5341 : STD_LOGIC;
    SIGNAL S5342 : STD_LOGIC;
    SIGNAL S5343 : STD_LOGIC;
    SIGNAL S5344 : STD_LOGIC;
    SIGNAL S5345 : STD_LOGIC;
    SIGNAL S5346 : STD_LOGIC;
    SIGNAL S5347 : STD_LOGIC;
    SIGNAL S5348 : STD_LOGIC;
    SIGNAL S5349 : STD_LOGIC;
    SIGNAL S5350 : STD_LOGIC;
    SIGNAL S5351 : STD_LOGIC;
    SIGNAL S5352 : STD_LOGIC;
    SIGNAL S5353 : STD_LOGIC;
    SIGNAL S5354 : STD_LOGIC;
    SIGNAL S5355 : STD_LOGIC;
    SIGNAL S5356 : STD_LOGIC;
    SIGNAL S5357 : STD_LOGIC;
    SIGNAL S5358 : STD_LOGIC;
    SIGNAL S5359 : STD_LOGIC;
    SIGNAL S5360 : STD_LOGIC;
    SIGNAL S5361 : STD_LOGIC;
    SIGNAL S5362 : STD_LOGIC;
    SIGNAL S5363 : STD_LOGIC;
    SIGNAL S5364 : STD_LOGIC;
    SIGNAL S5365 : STD_LOGIC;
    SIGNAL S5366 : STD_LOGIC;
    SIGNAL S5367 : STD_LOGIC;
    SIGNAL S5368 : STD_LOGIC;
    SIGNAL S5369 : STD_LOGIC;
    SIGNAL S5370 : STD_LOGIC;
    SIGNAL S5371 : STD_LOGIC;
    SIGNAL S5372 : STD_LOGIC;
    SIGNAL S5373 : STD_LOGIC;
    SIGNAL S5374 : STD_LOGIC;
    SIGNAL S5375 : STD_LOGIC;
    SIGNAL S5376 : STD_LOGIC;
    SIGNAL S5377 : STD_LOGIC;
    SIGNAL S5378 : STD_LOGIC;
    SIGNAL S5379 : STD_LOGIC;
    SIGNAL S5380 : STD_LOGIC;
    SIGNAL S5381 : STD_LOGIC;
    SIGNAL S5382 : STD_LOGIC;
    SIGNAL S5383 : STD_LOGIC;
    SIGNAL S5384 : STD_LOGIC;
    SIGNAL S5385 : STD_LOGIC;
    SIGNAL S5386 : STD_LOGIC;
    SIGNAL S5387 : STD_LOGIC;
    SIGNAL S5388 : STD_LOGIC;
    SIGNAL S5389 : STD_LOGIC;
    SIGNAL S5390 : STD_LOGIC;
    SIGNAL S5391 : STD_LOGIC;
    SIGNAL S5392 : STD_LOGIC;
    SIGNAL S5393 : STD_LOGIC;
    SIGNAL S5394 : STD_LOGIC;
    SIGNAL S5395 : STD_LOGIC;
    SIGNAL S5396 : STD_LOGIC;
    SIGNAL S5397 : STD_LOGIC;
    SIGNAL S5398 : STD_LOGIC;
    SIGNAL S5399 : STD_LOGIC;
    SIGNAL S5400 : STD_LOGIC;
    SIGNAL S5401 : STD_LOGIC;
    SIGNAL S5402 : STD_LOGIC;
    SIGNAL S5403 : STD_LOGIC;
    SIGNAL S5404 : STD_LOGIC;
    SIGNAL S5405 : STD_LOGIC;
    SIGNAL S5406 : STD_LOGIC;
    SIGNAL S5407 : STD_LOGIC;
    SIGNAL S5408 : STD_LOGIC;
    SIGNAL S5409 : STD_LOGIC;
    SIGNAL S5410 : STD_LOGIC;
    SIGNAL S5411 : STD_LOGIC;
    SIGNAL S5412 : STD_LOGIC;
    SIGNAL S5413 : STD_LOGIC;
    SIGNAL S5414 : STD_LOGIC;
    SIGNAL S5415 : STD_LOGIC;
    SIGNAL S5416 : STD_LOGIC;
    SIGNAL S5417 : STD_LOGIC;
    SIGNAL S5418 : STD_LOGIC;
    SIGNAL S5419 : STD_LOGIC;
    SIGNAL S5420 : STD_LOGIC;
    SIGNAL S5421 : STD_LOGIC;
    SIGNAL S5422 : STD_LOGIC;
    SIGNAL S5423 : STD_LOGIC;
    SIGNAL S5424 : STD_LOGIC;
    SIGNAL S5425 : STD_LOGIC;
    SIGNAL S5426 : STD_LOGIC;
    SIGNAL S5427 : STD_LOGIC;
    SIGNAL S5428 : STD_LOGIC;
    SIGNAL S5429 : STD_LOGIC;
    SIGNAL S5430 : STD_LOGIC;
    SIGNAL S5431 : STD_LOGIC;
    SIGNAL S5432 : STD_LOGIC;
    SIGNAL S5433 : STD_LOGIC;
    SIGNAL S5434 : STD_LOGIC;
    SIGNAL S5435 : STD_LOGIC;
    SIGNAL S5436 : STD_LOGIC;
    SIGNAL S5437 : STD_LOGIC;
    SIGNAL S5438 : STD_LOGIC;
    SIGNAL S5439 : STD_LOGIC;
    SIGNAL S5440 : STD_LOGIC;
    SIGNAL S5441 : STD_LOGIC;
    SIGNAL S5442 : STD_LOGIC;
    SIGNAL S5443 : STD_LOGIC;
    SIGNAL S5444 : STD_LOGIC;
    SIGNAL S5445 : STD_LOGIC;
    SIGNAL S5446 : STD_LOGIC;
    SIGNAL S5447 : STD_LOGIC;
    SIGNAL S5448 : STD_LOGIC;
    SIGNAL S5449 : STD_LOGIC;
    SIGNAL S5450 : STD_LOGIC;
    SIGNAL S5451 : STD_LOGIC;
    SIGNAL S5452 : STD_LOGIC;
    SIGNAL S5453 : STD_LOGIC;
    SIGNAL S5454 : STD_LOGIC;
    SIGNAL S5455 : STD_LOGIC;
    SIGNAL S5456 : STD_LOGIC;
    SIGNAL S5457 : STD_LOGIC;
    SIGNAL S5458 : STD_LOGIC;
    SIGNAL S5459 : STD_LOGIC;
    SIGNAL S5460 : STD_LOGIC;
    SIGNAL S5461 : STD_LOGIC;
    SIGNAL S5462 : STD_LOGIC;
    SIGNAL S5463 : STD_LOGIC;
    SIGNAL S5464 : STD_LOGIC;
    SIGNAL S5465 : STD_LOGIC;
    SIGNAL S5466 : STD_LOGIC;
    SIGNAL S5467 : STD_LOGIC;
    SIGNAL S5468 : STD_LOGIC;
    SIGNAL S5469 : STD_LOGIC;
    SIGNAL S5470 : STD_LOGIC;
    SIGNAL S5471 : STD_LOGIC;
    SIGNAL S5472 : STD_LOGIC;
    SIGNAL S5473 : STD_LOGIC;
    SIGNAL S5474 : STD_LOGIC;
    SIGNAL S5475 : STD_LOGIC;
    SIGNAL S5476 : STD_LOGIC;
    SIGNAL S5477 : STD_LOGIC;
    SIGNAL S5478 : STD_LOGIC;
    SIGNAL S5479 : STD_LOGIC;
    SIGNAL S5480 : STD_LOGIC;
    SIGNAL S5481 : STD_LOGIC;
    SIGNAL S5482 : STD_LOGIC;
    SIGNAL S5483 : STD_LOGIC;
    SIGNAL S5484 : STD_LOGIC;
    SIGNAL S5485 : STD_LOGIC;
    SIGNAL S5486 : STD_LOGIC;
    SIGNAL S5487 : STD_LOGIC;
    SIGNAL S5488 : STD_LOGIC;
    SIGNAL S5489 : STD_LOGIC;
    SIGNAL S5490 : STD_LOGIC;
    SIGNAL S5491 : STD_LOGIC;
    SIGNAL S5492 : STD_LOGIC;
    SIGNAL S5493 : STD_LOGIC;
    SIGNAL S5494 : STD_LOGIC;
    SIGNAL S5495 : STD_LOGIC;
    SIGNAL S5496 : STD_LOGIC;
    SIGNAL S5497 : STD_LOGIC;
    SIGNAL S5498 : STD_LOGIC;
    SIGNAL S5499 : STD_LOGIC;
    SIGNAL S5500 : STD_LOGIC;
    SIGNAL S5501 : STD_LOGIC;
    SIGNAL S5502 : STD_LOGIC;
    SIGNAL S5503 : STD_LOGIC;
    SIGNAL S5504 : STD_LOGIC;
    SIGNAL S5505 : STD_LOGIC;
    SIGNAL S5506 : STD_LOGIC;
    SIGNAL S5507 : STD_LOGIC;
    SIGNAL S5508 : STD_LOGIC;
    SIGNAL S5509 : STD_LOGIC;
    SIGNAL S5510 : STD_LOGIC;
    SIGNAL S5511 : STD_LOGIC;
    SIGNAL S5512 : STD_LOGIC;
    SIGNAL S5513 : STD_LOGIC;
    SIGNAL S5514 : STD_LOGIC;
    SIGNAL S5515 : STD_LOGIC;
    SIGNAL S5516 : STD_LOGIC;
    SIGNAL S5517 : STD_LOGIC;
    SIGNAL S5518 : STD_LOGIC;
    SIGNAL S5519 : STD_LOGIC;
    SIGNAL S5520 : STD_LOGIC;
    SIGNAL S5521 : STD_LOGIC;
    SIGNAL S5522 : STD_LOGIC;
    SIGNAL S5523 : STD_LOGIC;
    SIGNAL S5524 : STD_LOGIC;
    SIGNAL S5525 : STD_LOGIC;
    SIGNAL S5526 : STD_LOGIC;
    SIGNAL S5527 : STD_LOGIC;
    SIGNAL S5528 : STD_LOGIC;
    SIGNAL S5529 : STD_LOGIC;
    SIGNAL S5530 : STD_LOGIC;
    SIGNAL S5531 : STD_LOGIC;
    SIGNAL S5532 : STD_LOGIC;
    SIGNAL S5533 : STD_LOGIC;
    SIGNAL S5534 : STD_LOGIC;
    SIGNAL S5535 : STD_LOGIC;
    SIGNAL S5536 : STD_LOGIC;
    SIGNAL S5537 : STD_LOGIC;
    SIGNAL S5538 : STD_LOGIC;
    SIGNAL S5539 : STD_LOGIC;
    SIGNAL S5540 : STD_LOGIC;
    SIGNAL S5541 : STD_LOGIC;
    SIGNAL S5542 : STD_LOGIC;
    SIGNAL S5543 : STD_LOGIC;
    SIGNAL S5544 : STD_LOGIC;
    SIGNAL S5545 : STD_LOGIC;
    SIGNAL S5546 : STD_LOGIC;
    SIGNAL S5547 : STD_LOGIC;
    SIGNAL S5548 : STD_LOGIC;
    SIGNAL S5549 : STD_LOGIC;
    SIGNAL S5550 : STD_LOGIC;
    SIGNAL S5551 : STD_LOGIC;
    SIGNAL S5552 : STD_LOGIC;
    SIGNAL S5553 : STD_LOGIC;
    SIGNAL S5554 : STD_LOGIC;
    SIGNAL S5555 : STD_LOGIC;
    SIGNAL S5556 : STD_LOGIC;
    SIGNAL S5557 : STD_LOGIC;
    SIGNAL S5558 : STD_LOGIC;
    SIGNAL S5559 : STD_LOGIC;
    SIGNAL S5560 : STD_LOGIC;
    SIGNAL S5561 : STD_LOGIC;
    SIGNAL S5562 : STD_LOGIC;
    SIGNAL S5563 : STD_LOGIC;
    SIGNAL S5564 : STD_LOGIC;
    SIGNAL S5565 : STD_LOGIC;
    SIGNAL S5566 : STD_LOGIC;
    SIGNAL S5567 : STD_LOGIC;
    SIGNAL S5568 : STD_LOGIC;
    SIGNAL S5569 : STD_LOGIC;
    SIGNAL S5570 : STD_LOGIC;
    SIGNAL S5571 : STD_LOGIC;
    SIGNAL S5572 : STD_LOGIC;
    SIGNAL S5573 : STD_LOGIC;
    SIGNAL S5574 : STD_LOGIC;
    SIGNAL S5575 : STD_LOGIC;
    SIGNAL S5576 : STD_LOGIC;
    SIGNAL S5577 : STD_LOGIC;
    SIGNAL S5578 : STD_LOGIC;
    SIGNAL S5579 : STD_LOGIC;
    SIGNAL S5580 : STD_LOGIC;
    SIGNAL S5581 : STD_LOGIC;
    SIGNAL S5582 : STD_LOGIC;
    SIGNAL S5583 : STD_LOGIC;
    SIGNAL S5584 : STD_LOGIC;
    SIGNAL S5585 : STD_LOGIC;
    SIGNAL S5586 : STD_LOGIC;
    SIGNAL S5587 : STD_LOGIC;
    SIGNAL S5588 : STD_LOGIC;
    SIGNAL S5589 : STD_LOGIC;
    SIGNAL S5590 : STD_LOGIC;
    SIGNAL S5591 : STD_LOGIC;
    SIGNAL S5592 : STD_LOGIC;
    SIGNAL S5593 : STD_LOGIC;
    SIGNAL S5594 : STD_LOGIC;
    SIGNAL S5595 : STD_LOGIC;
    SIGNAL S5596 : STD_LOGIC;
    SIGNAL S5597 : STD_LOGIC;
    SIGNAL S5598 : STD_LOGIC;
    SIGNAL S5599 : STD_LOGIC;
    SIGNAL S5600 : STD_LOGIC;
    SIGNAL S5601 : STD_LOGIC;
    SIGNAL S5602 : STD_LOGIC;
    SIGNAL S5603 : STD_LOGIC;
    SIGNAL S5604 : STD_LOGIC;
    SIGNAL S5605 : STD_LOGIC;
    SIGNAL S5606 : STD_LOGIC;
    SIGNAL S5607 : STD_LOGIC;
    SIGNAL S5608 : STD_LOGIC;
    SIGNAL S5609 : STD_LOGIC;
    SIGNAL S5610 : STD_LOGIC;
    SIGNAL S5611 : STD_LOGIC;
    SIGNAL S5612 : STD_LOGIC;
    SIGNAL S5613 : STD_LOGIC;
    SIGNAL S5614 : STD_LOGIC;
    SIGNAL S5615 : STD_LOGIC;
    SIGNAL S5616 : STD_LOGIC;
    SIGNAL S5617 : STD_LOGIC;
    SIGNAL S5618 : STD_LOGIC;
    SIGNAL S5619 : STD_LOGIC;
    SIGNAL S5620 : STD_LOGIC;
    SIGNAL S5621 : STD_LOGIC;
    SIGNAL S5622 : STD_LOGIC;
    SIGNAL S5623 : STD_LOGIC;
    SIGNAL S5624 : STD_LOGIC;
    SIGNAL S5625 : STD_LOGIC;
    SIGNAL S5626 : STD_LOGIC;
    SIGNAL S5627 : STD_LOGIC;
    SIGNAL S5628 : STD_LOGIC;
    SIGNAL S5629 : STD_LOGIC;
    SIGNAL S5630 : STD_LOGIC;
    SIGNAL S5631 : STD_LOGIC;
    SIGNAL S5632 : STD_LOGIC;
    SIGNAL S5633 : STD_LOGIC;
    SIGNAL S5634 : STD_LOGIC;
    SIGNAL S5635 : STD_LOGIC;
    SIGNAL S5636 : STD_LOGIC;
    SIGNAL S5637 : STD_LOGIC;
    SIGNAL S5638 : STD_LOGIC;
    SIGNAL S5639 : STD_LOGIC;
    SIGNAL S5640 : STD_LOGIC;
    SIGNAL S5641 : STD_LOGIC;
    SIGNAL S5642 : STD_LOGIC;
    SIGNAL S5643 : STD_LOGIC;
    SIGNAL S5644 : STD_LOGIC;
    SIGNAL S5645 : STD_LOGIC;
    SIGNAL S5646 : STD_LOGIC;
    SIGNAL S5647 : STD_LOGIC;
    SIGNAL S5648 : STD_LOGIC;
    SIGNAL S5649 : STD_LOGIC;
    SIGNAL S5650 : STD_LOGIC;
    SIGNAL S5651 : STD_LOGIC;
    SIGNAL S5652 : STD_LOGIC;
    SIGNAL S5653 : STD_LOGIC;
    SIGNAL S5654 : STD_LOGIC;
    SIGNAL S5655 : STD_LOGIC;
    SIGNAL S5656 : STD_LOGIC;
    SIGNAL S5657 : STD_LOGIC;
    SIGNAL S5658 : STD_LOGIC;
    SIGNAL S5659 : STD_LOGIC;
    SIGNAL S5660 : STD_LOGIC;
    SIGNAL S5661 : STD_LOGIC;
    SIGNAL S5662 : STD_LOGIC;
    SIGNAL S5663 : STD_LOGIC;
    SIGNAL S5664 : STD_LOGIC;
    SIGNAL S5665 : STD_LOGIC;
    SIGNAL S5666 : STD_LOGIC;
    SIGNAL S5667 : STD_LOGIC;
    SIGNAL S5668 : STD_LOGIC;
    SIGNAL S5669 : STD_LOGIC;
    SIGNAL S5670 : STD_LOGIC;
    SIGNAL S5671 : STD_LOGIC;
    SIGNAL S5672 : STD_LOGIC;
    SIGNAL S5673 : STD_LOGIC;
    SIGNAL S5674 : STD_LOGIC;
    SIGNAL S5675 : STD_LOGIC;
    SIGNAL S5676 : STD_LOGIC;
    SIGNAL S5677 : STD_LOGIC;
    SIGNAL S5678 : STD_LOGIC;
    SIGNAL S5679 : STD_LOGIC;
    SIGNAL S5680 : STD_LOGIC;
    SIGNAL S5681 : STD_LOGIC;
    SIGNAL S5682 : STD_LOGIC;
    SIGNAL S5683 : STD_LOGIC;
    SIGNAL S5684 : STD_LOGIC;
    SIGNAL S5685 : STD_LOGIC;
    SIGNAL S5686 : STD_LOGIC;
    SIGNAL S5687 : STD_LOGIC;
    SIGNAL S5688 : STD_LOGIC;
    SIGNAL S5689 : STD_LOGIC;
    SIGNAL S5690 : STD_LOGIC;
    SIGNAL S5691 : STD_LOGIC;
    SIGNAL S5692 : STD_LOGIC;
    SIGNAL S5693 : STD_LOGIC;
    SIGNAL S5694 : STD_LOGIC;
    SIGNAL S5695 : STD_LOGIC;
    SIGNAL S5696 : STD_LOGIC;
    SIGNAL S5697 : STD_LOGIC;
    SIGNAL S5698 : STD_LOGIC;
    SIGNAL S5699 : STD_LOGIC;
    SIGNAL S5700 : STD_LOGIC;
    SIGNAL S5701 : STD_LOGIC;
    SIGNAL S5702 : STD_LOGIC;
    SIGNAL S5703 : STD_LOGIC;
    SIGNAL S5704 : STD_LOGIC;
    SIGNAL S5705 : STD_LOGIC;
    SIGNAL S5706 : STD_LOGIC;
    SIGNAL S5707 : STD_LOGIC;
    SIGNAL S5708 : STD_LOGIC;
    SIGNAL S5709 : STD_LOGIC;
    SIGNAL S5710 : STD_LOGIC;
    SIGNAL S5711 : STD_LOGIC;
    SIGNAL S5712 : STD_LOGIC;
    SIGNAL S5713 : STD_LOGIC;
    SIGNAL S5714 : STD_LOGIC;
    SIGNAL S5715 : STD_LOGIC;
    SIGNAL S5716 : STD_LOGIC;
    SIGNAL S5717 : STD_LOGIC;
    SIGNAL S5718 : STD_LOGIC;
    SIGNAL S5719 : STD_LOGIC;
    SIGNAL S5720 : STD_LOGIC;
    SIGNAL S5721 : STD_LOGIC;
    SIGNAL S5722 : STD_LOGIC;
    SIGNAL S5723 : STD_LOGIC;
    SIGNAL S5724 : STD_LOGIC;
    SIGNAL S5725 : STD_LOGIC;
    SIGNAL S5726 : STD_LOGIC;
    SIGNAL S5727 : STD_LOGIC;
    SIGNAL S5728 : STD_LOGIC;
    SIGNAL S5729 : STD_LOGIC;
    SIGNAL S5730 : STD_LOGIC;
    SIGNAL S5731 : STD_LOGIC;
    SIGNAL S5732 : STD_LOGIC;
    SIGNAL S5733 : STD_LOGIC;
    SIGNAL S5734 : STD_LOGIC;
    SIGNAL S5735 : STD_LOGIC;
    SIGNAL S5736 : STD_LOGIC;
    SIGNAL S5737 : STD_LOGIC;
    SIGNAL S5738 : STD_LOGIC;
    SIGNAL S5739 : STD_LOGIC;
    SIGNAL S5740 : STD_LOGIC;
    SIGNAL S5741 : STD_LOGIC;
    SIGNAL S5742 : STD_LOGIC;
    SIGNAL S5743 : STD_LOGIC;
    SIGNAL S5744 : STD_LOGIC;
    SIGNAL S5745 : STD_LOGIC;
    SIGNAL S5746 : STD_LOGIC;
    SIGNAL S5747 : STD_LOGIC;
    SIGNAL S5748 : STD_LOGIC;
    SIGNAL S5749 : STD_LOGIC;
    SIGNAL S5750 : STD_LOGIC;
    SIGNAL S5751 : STD_LOGIC;
    SIGNAL S5752 : STD_LOGIC;
    SIGNAL S5753 : STD_LOGIC;
    SIGNAL S5754 : STD_LOGIC;
    SIGNAL S5755 : STD_LOGIC;
    SIGNAL S5756 : STD_LOGIC;
    SIGNAL S5757 : STD_LOGIC;
    SIGNAL S5758 : STD_LOGIC;
    SIGNAL S5759 : STD_LOGIC;
    SIGNAL S5760 : STD_LOGIC;
    SIGNAL S5761 : STD_LOGIC;
    SIGNAL S5762 : STD_LOGIC;
    SIGNAL S5763 : STD_LOGIC;
    SIGNAL S5764 : STD_LOGIC;
    SIGNAL S5765 : STD_LOGIC;
    SIGNAL S5766 : STD_LOGIC;
    SIGNAL S5767 : STD_LOGIC;
    SIGNAL S5768 : STD_LOGIC;
    SIGNAL S5769 : STD_LOGIC;
    SIGNAL S5770 : STD_LOGIC;
    SIGNAL S5771 : STD_LOGIC;
    SIGNAL S5772 : STD_LOGIC;
    SIGNAL S5773 : STD_LOGIC;
    SIGNAL S5774 : STD_LOGIC;
    SIGNAL S5775 : STD_LOGIC;
    SIGNAL S5776 : STD_LOGIC;
    SIGNAL S5777 : STD_LOGIC;
    SIGNAL S5778 : STD_LOGIC;
    SIGNAL S5779 : STD_LOGIC;
    SIGNAL S5780 : STD_LOGIC;
    SIGNAL S5781 : STD_LOGIC;
    SIGNAL S5782 : STD_LOGIC;
    SIGNAL S5783 : STD_LOGIC;
    SIGNAL S5784 : STD_LOGIC;
    SIGNAL S5785 : STD_LOGIC;
    SIGNAL S5786 : STD_LOGIC;
    SIGNAL S5787 : STD_LOGIC;
    SIGNAL S5788 : STD_LOGIC;
    SIGNAL S5789 : STD_LOGIC;
    SIGNAL S5790 : STD_LOGIC;
    SIGNAL S5791 : STD_LOGIC;
    SIGNAL S5792 : STD_LOGIC;
    SIGNAL S5793 : STD_LOGIC;
    SIGNAL S5794 : STD_LOGIC;
    SIGNAL S5795 : STD_LOGIC;
    SIGNAL S5796 : STD_LOGIC;
    SIGNAL S5797 : STD_LOGIC;
    SIGNAL S5798 : STD_LOGIC;
    SIGNAL S5799 : STD_LOGIC;
    SIGNAL S5800 : STD_LOGIC;
    SIGNAL S5801 : STD_LOGIC;
    SIGNAL S5802 : STD_LOGIC;
    SIGNAL S5803 : STD_LOGIC;
    SIGNAL S5804 : STD_LOGIC;
    SIGNAL S5805 : STD_LOGIC;
    SIGNAL S5806 : STD_LOGIC;
    SIGNAL S5807 : STD_LOGIC;
    SIGNAL S5808 : STD_LOGIC;
    SIGNAL S5809 : STD_LOGIC;
    SIGNAL S5810 : STD_LOGIC;
    SIGNAL S5811 : STD_LOGIC;
    SIGNAL S5812 : STD_LOGIC;
    SIGNAL S5813 : STD_LOGIC;
    SIGNAL S5814 : STD_LOGIC;
    SIGNAL S5815 : STD_LOGIC;
    SIGNAL S5816 : STD_LOGIC;
    SIGNAL S5817 : STD_LOGIC;
    SIGNAL S5818 : STD_LOGIC;
    SIGNAL S5819 : STD_LOGIC;
    SIGNAL S5820 : STD_LOGIC;
    SIGNAL S5821 : STD_LOGIC;
    SIGNAL S5822 : STD_LOGIC;
    SIGNAL S5823 : STD_LOGIC;
    SIGNAL S5824 : STD_LOGIC;
    SIGNAL S5825 : STD_LOGIC;
    SIGNAL S5826 : STD_LOGIC;
    SIGNAL S5827 : STD_LOGIC;
    SIGNAL S5828 : STD_LOGIC;
    SIGNAL S5829 : STD_LOGIC;
    SIGNAL S5830 : STD_LOGIC;
    SIGNAL S5831 : STD_LOGIC;
    SIGNAL S5832 : STD_LOGIC;
    SIGNAL S5833 : STD_LOGIC;
    SIGNAL S5834 : STD_LOGIC;
    SIGNAL S5835 : STD_LOGIC;
    SIGNAL S5836 : STD_LOGIC;
    SIGNAL S5837 : STD_LOGIC;
    SIGNAL S5838 : STD_LOGIC;
    SIGNAL S5839 : STD_LOGIC;
    SIGNAL S5840 : STD_LOGIC;
    SIGNAL S5841 : STD_LOGIC;
    SIGNAL S5842 : STD_LOGIC;
    SIGNAL S5843 : STD_LOGIC;
    SIGNAL S5844 : STD_LOGIC;
    SIGNAL S5845 : STD_LOGIC;
    SIGNAL S5846 : STD_LOGIC;
    SIGNAL S5847 : STD_LOGIC;
    SIGNAL S5848 : STD_LOGIC;
    SIGNAL S5849 : STD_LOGIC;
    SIGNAL S5850 : STD_LOGIC;
    SIGNAL S5851 : STD_LOGIC;
    SIGNAL S5852 : STD_LOGIC;
    SIGNAL S5853 : STD_LOGIC;
    SIGNAL S5854 : STD_LOGIC;
    SIGNAL S5855 : STD_LOGIC;
    SIGNAL S5856 : STD_LOGIC;
    SIGNAL S5857 : STD_LOGIC;
    SIGNAL S5858 : STD_LOGIC;
    SIGNAL S5859 : STD_LOGIC;
    SIGNAL S5860 : STD_LOGIC;
    SIGNAL S5861 : STD_LOGIC;
    SIGNAL S5862 : STD_LOGIC;
    SIGNAL S5863 : STD_LOGIC;
    SIGNAL S5864 : STD_LOGIC;
    SIGNAL S5865 : STD_LOGIC;
    SIGNAL S5866 : STD_LOGIC;
    SIGNAL S5867 : STD_LOGIC;
    SIGNAL S5868 : STD_LOGIC;
    SIGNAL S5869 : STD_LOGIC;
    SIGNAL S5870 : STD_LOGIC;
    SIGNAL S5871 : STD_LOGIC;
    SIGNAL S5872 : STD_LOGIC;
    SIGNAL S5873 : STD_LOGIC;
    SIGNAL S5874 : STD_LOGIC;
    SIGNAL S5875 : STD_LOGIC;
    SIGNAL S5876 : STD_LOGIC;
    SIGNAL S5877 : STD_LOGIC;
    SIGNAL S5878 : STD_LOGIC;
    SIGNAL S5879 : STD_LOGIC;
    SIGNAL S5880 : STD_LOGIC;
    SIGNAL S5881 : STD_LOGIC;
    SIGNAL S5882 : STD_LOGIC;
    SIGNAL S5883 : STD_LOGIC;
    SIGNAL S5884 : STD_LOGIC;
    SIGNAL S5885 : STD_LOGIC;
    SIGNAL S5886 : STD_LOGIC;
    SIGNAL S5887 : STD_LOGIC;
    SIGNAL S5888 : STD_LOGIC;
    SIGNAL S5889 : STD_LOGIC;
    SIGNAL S5890 : STD_LOGIC;
    SIGNAL S5891 : STD_LOGIC;
    SIGNAL S5892 : STD_LOGIC;
    SIGNAL S5893 : STD_LOGIC;
    SIGNAL S5894 : STD_LOGIC;
    SIGNAL S5895 : STD_LOGIC;
    SIGNAL S5896 : STD_LOGIC;
    SIGNAL S5897 : STD_LOGIC;
    SIGNAL S5898 : STD_LOGIC;
    SIGNAL S5899 : STD_LOGIC;
    SIGNAL S5900 : STD_LOGIC;
    SIGNAL S5901 : STD_LOGIC;
    SIGNAL S5902 : STD_LOGIC;
    SIGNAL S5903 : STD_LOGIC;
    SIGNAL S5904 : STD_LOGIC;
    SIGNAL S5905 : STD_LOGIC;
    SIGNAL S5906 : STD_LOGIC;
    SIGNAL S5907 : STD_LOGIC;
    SIGNAL S5908 : STD_LOGIC;
    SIGNAL S5909 : STD_LOGIC;
    SIGNAL S5910 : STD_LOGIC;
    SIGNAL S5911 : STD_LOGIC;
    SIGNAL S5912 : STD_LOGIC;
    SIGNAL S5913 : STD_LOGIC;
    SIGNAL S5914 : STD_LOGIC;
    SIGNAL S5915 : STD_LOGIC;
    SIGNAL S5916 : STD_LOGIC;
    SIGNAL S5917 : STD_LOGIC;
    SIGNAL S5918 : STD_LOGIC;
    SIGNAL S5919 : STD_LOGIC;
    SIGNAL S5920 : STD_LOGIC;
    SIGNAL S5921 : STD_LOGIC;
    SIGNAL S5922 : STD_LOGIC;
    SIGNAL S5923 : STD_LOGIC;
    SIGNAL S5924 : STD_LOGIC;
    SIGNAL S5925 : STD_LOGIC;
    SIGNAL S5926 : STD_LOGIC;
    SIGNAL S5927 : STD_LOGIC;
    SIGNAL S5928 : STD_LOGIC;
    SIGNAL S5929 : STD_LOGIC;
    SIGNAL S5930 : STD_LOGIC;
    SIGNAL S5931 : STD_LOGIC;
    SIGNAL S5932 : STD_LOGIC;
    SIGNAL S5933 : STD_LOGIC;
    SIGNAL S5934 : STD_LOGIC;
    SIGNAL S5935 : STD_LOGIC;
    SIGNAL S5936 : STD_LOGIC;
    SIGNAL S5937 : STD_LOGIC;
    SIGNAL S5938 : STD_LOGIC;
    SIGNAL S5939 : STD_LOGIC;
    SIGNAL S5940 : STD_LOGIC;
    SIGNAL S5941 : STD_LOGIC;
    SIGNAL S5942 : STD_LOGIC;
    SIGNAL S5943 : STD_LOGIC;
    SIGNAL S5944 : STD_LOGIC;
    SIGNAL S5945 : STD_LOGIC;
    SIGNAL S5946 : STD_LOGIC;
    SIGNAL S5947 : STD_LOGIC;
    SIGNAL S5948 : STD_LOGIC;
    SIGNAL S5949 : STD_LOGIC;
    SIGNAL S5950 : STD_LOGIC;
    SIGNAL S5951 : STD_LOGIC;
    SIGNAL S5952 : STD_LOGIC;
    SIGNAL S5953 : STD_LOGIC;
    SIGNAL S5954 : STD_LOGIC;
    SIGNAL S5955 : STD_LOGIC;
    SIGNAL S5956 : STD_LOGIC;
    SIGNAL S5957 : STD_LOGIC;
    SIGNAL S5958 : STD_LOGIC;
    SIGNAL S5959 : STD_LOGIC;
    SIGNAL S5960 : STD_LOGIC;
    SIGNAL S5961 : STD_LOGIC;
    SIGNAL S5962 : STD_LOGIC;
    SIGNAL S5963 : STD_LOGIC;
    SIGNAL S5964 : STD_LOGIC;
    SIGNAL S5965 : STD_LOGIC;
    SIGNAL S5966 : STD_LOGIC;
    SIGNAL S5967 : STD_LOGIC;
    SIGNAL S5968 : STD_LOGIC;
    SIGNAL S5969 : STD_LOGIC;
    SIGNAL S5970 : STD_LOGIC;
    SIGNAL S5971 : STD_LOGIC;
    SIGNAL S5972 : STD_LOGIC;
    SIGNAL S5973 : STD_LOGIC;
    SIGNAL S5974 : STD_LOGIC;
    SIGNAL S5975 : STD_LOGIC;
    SIGNAL S5976 : STD_LOGIC;
    SIGNAL S5977 : STD_LOGIC;
    SIGNAL S5978 : STD_LOGIC;
    SIGNAL S5979 : STD_LOGIC;
    SIGNAL S5980 : STD_LOGIC;
    SIGNAL S5981 : STD_LOGIC;
    SIGNAL S5982 : STD_LOGIC;
    SIGNAL S5983 : STD_LOGIC;
    SIGNAL S5984 : STD_LOGIC;
    SIGNAL S5985 : STD_LOGIC;
    SIGNAL S5986 : STD_LOGIC;
    SIGNAL S5987 : STD_LOGIC;
    SIGNAL S5988 : STD_LOGIC;
    SIGNAL S5989 : STD_LOGIC;
    SIGNAL S5990 : STD_LOGIC;
    SIGNAL S5991 : STD_LOGIC;
    SIGNAL S5992 : STD_LOGIC;
    SIGNAL S5993 : STD_LOGIC;
    SIGNAL S5994 : STD_LOGIC;
    SIGNAL S5995 : STD_LOGIC;
    SIGNAL S5996 : STD_LOGIC;
    SIGNAL S5997 : STD_LOGIC;
    SIGNAL S5998 : STD_LOGIC;
    SIGNAL S5999 : STD_LOGIC;
    SIGNAL S6000 : STD_LOGIC;
    SIGNAL S6001 : STD_LOGIC;
    SIGNAL S6002 : STD_LOGIC;
    SIGNAL S6003 : STD_LOGIC;
    SIGNAL S6004 : STD_LOGIC;
    SIGNAL S6005 : STD_LOGIC;
    SIGNAL S6006 : STD_LOGIC;
    SIGNAL S6007 : STD_LOGIC;
    SIGNAL S6008 : STD_LOGIC;
    SIGNAL S6009 : STD_LOGIC;
    SIGNAL S6010 : STD_LOGIC;
    SIGNAL S6011 : STD_LOGIC;
    SIGNAL S6012 : STD_LOGIC;
    SIGNAL S6013 : STD_LOGIC;
    SIGNAL S6014 : STD_LOGIC;
    SIGNAL S6015 : STD_LOGIC;
    SIGNAL S6016 : STD_LOGIC;
    SIGNAL S6017 : STD_LOGIC;
    SIGNAL S6018 : STD_LOGIC;
    SIGNAL S6019 : STD_LOGIC;
    SIGNAL S6020 : STD_LOGIC;
    SIGNAL S6021 : STD_LOGIC;
    SIGNAL S6022 : STD_LOGIC;
    SIGNAL S6023 : STD_LOGIC;
    SIGNAL S6024 : STD_LOGIC;
    SIGNAL S6025 : STD_LOGIC;
    SIGNAL S6026 : STD_LOGIC;
    SIGNAL S6027 : STD_LOGIC;
    SIGNAL S6028 : STD_LOGIC;
    SIGNAL S6029 : STD_LOGIC;
    SIGNAL S6030 : STD_LOGIC;
    SIGNAL S6031 : STD_LOGIC;
    SIGNAL S6032 : STD_LOGIC;
    SIGNAL S6033 : STD_LOGIC;
    SIGNAL S6034 : STD_LOGIC;
    SIGNAL S6035 : STD_LOGIC;
    SIGNAL S6036 : STD_LOGIC;
    SIGNAL S6037 : STD_LOGIC;
    SIGNAL S6038 : STD_LOGIC;
    SIGNAL S6039 : STD_LOGIC;
    SIGNAL S6040 : STD_LOGIC;
    SIGNAL S6041 : STD_LOGIC;
    SIGNAL S6042 : STD_LOGIC;
    SIGNAL S6043 : STD_LOGIC;
    SIGNAL S6044 : STD_LOGIC;
    SIGNAL S6045 : STD_LOGIC;
    SIGNAL S6046 : STD_LOGIC;
    SIGNAL S6047 : STD_LOGIC;
    SIGNAL S6048 : STD_LOGIC;
    SIGNAL S6049 : STD_LOGIC;
    SIGNAL S6050 : STD_LOGIC;
    SIGNAL S6051 : STD_LOGIC;
    SIGNAL S6052 : STD_LOGIC;
    SIGNAL S6053 : STD_LOGIC;
    SIGNAL S6054 : STD_LOGIC;
    SIGNAL S6055 : STD_LOGIC;
    SIGNAL S6056 : STD_LOGIC;
    SIGNAL S6057 : STD_LOGIC;
    SIGNAL S6058 : STD_LOGIC;
    SIGNAL S6059 : STD_LOGIC;
    SIGNAL S6060 : STD_LOGIC;
    SIGNAL S6061 : STD_LOGIC;
    SIGNAL S6062 : STD_LOGIC;
    SIGNAL S6063 : STD_LOGIC;
    SIGNAL S6064 : STD_LOGIC;
    SIGNAL S6065 : STD_LOGIC;
    SIGNAL S6066 : STD_LOGIC;
    SIGNAL S6067 : STD_LOGIC;
    SIGNAL S6068 : STD_LOGIC;
    SIGNAL S6069 : STD_LOGIC;
    SIGNAL S6070 : STD_LOGIC;
    SIGNAL S6071 : STD_LOGIC;
    SIGNAL S6072 : STD_LOGIC;
    SIGNAL S6073 : STD_LOGIC;
    SIGNAL S6074 : STD_LOGIC;
    SIGNAL S6075 : STD_LOGIC;
    SIGNAL S6076 : STD_LOGIC;
    SIGNAL S6077 : STD_LOGIC;
    SIGNAL S6078 : STD_LOGIC;
    SIGNAL S6079 : STD_LOGIC;
    SIGNAL S6080 : STD_LOGIC;
    SIGNAL S6081 : STD_LOGIC;
    SIGNAL S6082 : STD_LOGIC;
    SIGNAL S6083 : STD_LOGIC;
    SIGNAL S6084 : STD_LOGIC;
    SIGNAL S6085 : STD_LOGIC;
    SIGNAL S6086 : STD_LOGIC;
    SIGNAL S6087 : STD_LOGIC;
    SIGNAL S6088 : STD_LOGIC;
    SIGNAL S6089 : STD_LOGIC;
    SIGNAL S6090 : STD_LOGIC;
    SIGNAL S6091 : STD_LOGIC;
    SIGNAL S6092 : STD_LOGIC;
    SIGNAL S6093 : STD_LOGIC;
    SIGNAL S6094 : STD_LOGIC;
    SIGNAL S6095 : STD_LOGIC;
    SIGNAL S6096 : STD_LOGIC;
    SIGNAL S6097 : STD_LOGIC;
    SIGNAL S6098 : STD_LOGIC;
    SIGNAL S6099 : STD_LOGIC;
    SIGNAL S6100 : STD_LOGIC;
    SIGNAL S6101 : STD_LOGIC;
    SIGNAL S6102 : STD_LOGIC;
    SIGNAL S6103 : STD_LOGIC;
    SIGNAL S6104 : STD_LOGIC;
    SIGNAL S6105 : STD_LOGIC;
    SIGNAL S6106 : STD_LOGIC;
    SIGNAL S6107 : STD_LOGIC;
    SIGNAL S6108 : STD_LOGIC;
    SIGNAL S6109 : STD_LOGIC;
    SIGNAL S6110 : STD_LOGIC;
    SIGNAL S6111 : STD_LOGIC;
    SIGNAL S6112 : STD_LOGIC;
    SIGNAL S6113 : STD_LOGIC;
    SIGNAL S6114 : STD_LOGIC;
    SIGNAL S6115 : STD_LOGIC;
    SIGNAL S6116 : STD_LOGIC;
    SIGNAL S6117 : STD_LOGIC;
    SIGNAL S6118 : STD_LOGIC;
    SIGNAL S6119 : STD_LOGIC;
    SIGNAL S6120 : STD_LOGIC;
    SIGNAL S6121 : STD_LOGIC;
    SIGNAL S6122 : STD_LOGIC;
    SIGNAL S6123 : STD_LOGIC;
    SIGNAL S6124 : STD_LOGIC;
    SIGNAL S6125 : STD_LOGIC;
    SIGNAL S6126 : STD_LOGIC;
    SIGNAL S6127 : STD_LOGIC;
    SIGNAL S6128 : STD_LOGIC;
    SIGNAL S6129 : STD_LOGIC;
    SIGNAL S6130 : STD_LOGIC;
    SIGNAL S6131 : STD_LOGIC;
    SIGNAL S6132 : STD_LOGIC;
    SIGNAL S6133 : STD_LOGIC;
    SIGNAL S6134 : STD_LOGIC;
    SIGNAL S6135 : STD_LOGIC;
    SIGNAL S6136 : STD_LOGIC;
    SIGNAL S6137 : STD_LOGIC;
    SIGNAL S6138 : STD_LOGIC;
    SIGNAL S6139 : STD_LOGIC;
    SIGNAL S6140 : STD_LOGIC;
    SIGNAL S6141 : STD_LOGIC;
    SIGNAL S6142 : STD_LOGIC;
    SIGNAL S6143 : STD_LOGIC;
    SIGNAL S6144 : STD_LOGIC;
    SIGNAL S6145 : STD_LOGIC;
    SIGNAL S6146 : STD_LOGIC;
    SIGNAL S6147 : STD_LOGIC;
    SIGNAL S6148 : STD_LOGIC;
    SIGNAL S6149 : STD_LOGIC;
    SIGNAL S6150 : STD_LOGIC;
    SIGNAL S6151 : STD_LOGIC;
    SIGNAL S6152 : STD_LOGIC;
    SIGNAL S6153 : STD_LOGIC;
    SIGNAL S6154 : STD_LOGIC;
    SIGNAL S6155 : STD_LOGIC;
    SIGNAL S6156 : STD_LOGIC;
    SIGNAL S6157 : STD_LOGIC;
    SIGNAL S6158 : STD_LOGIC;
    SIGNAL S6159 : STD_LOGIC;
    SIGNAL S6160 : STD_LOGIC;
    SIGNAL S6161 : STD_LOGIC;
    SIGNAL S6162 : STD_LOGIC;
    SIGNAL S6163 : STD_LOGIC;
    SIGNAL S6164 : STD_LOGIC;
    SIGNAL S6165 : STD_LOGIC;
    SIGNAL S6166 : STD_LOGIC;
    SIGNAL S6167 : STD_LOGIC;
    SIGNAL S6168 : STD_LOGIC;
    SIGNAL S6169 : STD_LOGIC;
    SIGNAL S6170 : STD_LOGIC;
    SIGNAL S6171 : STD_LOGIC;
    SIGNAL S6172 : STD_LOGIC;
    SIGNAL S6173 : STD_LOGIC;
    SIGNAL S6174 : STD_LOGIC;
    SIGNAL S6175 : STD_LOGIC;
    SIGNAL S6176 : STD_LOGIC;
    SIGNAL S6177 : STD_LOGIC;
    SIGNAL S6178 : STD_LOGIC;
    SIGNAL S6179 : STD_LOGIC;
    SIGNAL S6180 : STD_LOGIC;
    SIGNAL S6181 : STD_LOGIC;
    SIGNAL S6182 : STD_LOGIC;
    SIGNAL S6183 : STD_LOGIC;
    SIGNAL S6184 : STD_LOGIC;
    SIGNAL S6185 : STD_LOGIC;
    SIGNAL S6186 : STD_LOGIC;
    SIGNAL S6187 : STD_LOGIC;
    SIGNAL S6188 : STD_LOGIC;
    SIGNAL S6189 : STD_LOGIC;
    SIGNAL S6190 : STD_LOGIC;
    SIGNAL S6191 : STD_LOGIC;
    SIGNAL S6192 : STD_LOGIC;
    SIGNAL S6193 : STD_LOGIC;
    SIGNAL S6194 : STD_LOGIC;
    SIGNAL S6195 : STD_LOGIC;
    SIGNAL S6196 : STD_LOGIC;
    SIGNAL S6197 : STD_LOGIC;
    SIGNAL S6198 : STD_LOGIC;
    SIGNAL S6199 : STD_LOGIC;
    SIGNAL S6200 : STD_LOGIC;
    SIGNAL S6201 : STD_LOGIC;
    SIGNAL S6202 : STD_LOGIC;
    SIGNAL S6203 : STD_LOGIC;
    SIGNAL S6204 : STD_LOGIC;
    SIGNAL S6205 : STD_LOGIC;
    SIGNAL S6206 : STD_LOGIC;
    SIGNAL S6207 : STD_LOGIC;
    SIGNAL S6208 : STD_LOGIC;
    SIGNAL S6209 : STD_LOGIC;
    SIGNAL S6210 : STD_LOGIC;
    SIGNAL S6211 : STD_LOGIC;
    SIGNAL S6212 : STD_LOGIC;
    SIGNAL S6213 : STD_LOGIC;
    SIGNAL S6214 : STD_LOGIC;
    SIGNAL S6215 : STD_LOGIC;
    SIGNAL S6216 : STD_LOGIC;
    SIGNAL S6217 : STD_LOGIC;
    SIGNAL S6218 : STD_LOGIC;
    SIGNAL S6219 : STD_LOGIC;
    SIGNAL S6220 : STD_LOGIC;
    SIGNAL S6221 : STD_LOGIC;
    SIGNAL S6222 : STD_LOGIC;
    SIGNAL S6223 : STD_LOGIC;
    SIGNAL S6224 : STD_LOGIC;
    SIGNAL S6225 : STD_LOGIC;
    SIGNAL S6226 : STD_LOGIC;
    SIGNAL S6227 : STD_LOGIC;
    SIGNAL S6228 : STD_LOGIC;
    SIGNAL S6229 : STD_LOGIC;
    SIGNAL S6230 : STD_LOGIC;
    SIGNAL S6231 : STD_LOGIC;
    SIGNAL S6232 : STD_LOGIC;
    SIGNAL S6233 : STD_LOGIC;
    SIGNAL S6234 : STD_LOGIC;
    SIGNAL S6235 : STD_LOGIC;
    SIGNAL S6236 : STD_LOGIC;
    SIGNAL S6237 : STD_LOGIC;
    SIGNAL S6238 : STD_LOGIC;
    SIGNAL S6239 : STD_LOGIC;
    SIGNAL S6240 : STD_LOGIC;
    SIGNAL S6241 : STD_LOGIC;
    SIGNAL S6242 : STD_LOGIC;
    SIGNAL S6243 : STD_LOGIC;
    SIGNAL S6244 : STD_LOGIC;
    SIGNAL S6245 : STD_LOGIC;
    SIGNAL S6246 : STD_LOGIC;
    SIGNAL S6247 : STD_LOGIC;
    SIGNAL S6248 : STD_LOGIC;
    SIGNAL S6249 : STD_LOGIC;
    SIGNAL S6250 : STD_LOGIC;
    SIGNAL S6251 : STD_LOGIC;
    SIGNAL S6252 : STD_LOGIC;
    SIGNAL S6253 : STD_LOGIC;
    SIGNAL S6254 : STD_LOGIC;
    SIGNAL S6255 : STD_LOGIC;
    SIGNAL S6256 : STD_LOGIC;
    SIGNAL S6257 : STD_LOGIC;
    SIGNAL S6258 : STD_LOGIC;
    SIGNAL S6259 : STD_LOGIC;
    SIGNAL S6260 : STD_LOGIC;
    SIGNAL S6261 : STD_LOGIC;
    SIGNAL S6262 : STD_LOGIC;
    SIGNAL S6263 : STD_LOGIC;
    SIGNAL S6264 : STD_LOGIC;
    SIGNAL S6265 : STD_LOGIC;
    SIGNAL S6266 : STD_LOGIC;
    SIGNAL S6267 : STD_LOGIC;
    SIGNAL S6268 : STD_LOGIC;
    SIGNAL S6269 : STD_LOGIC;
    SIGNAL S6270 : STD_LOGIC;
    SIGNAL S6271 : STD_LOGIC;
    SIGNAL S6272 : STD_LOGIC;
    SIGNAL S6273 : STD_LOGIC;
    SIGNAL S6274 : STD_LOGIC;
    SIGNAL S6275 : STD_LOGIC;
    SIGNAL S6276 : STD_LOGIC;
    SIGNAL S6277 : STD_LOGIC;
    SIGNAL S6278 : STD_LOGIC;
    SIGNAL S6279 : STD_LOGIC;
    SIGNAL S6280 : STD_LOGIC;
    SIGNAL S6281 : STD_LOGIC;
    SIGNAL S6282 : STD_LOGIC;
    SIGNAL S6283 : STD_LOGIC;
    SIGNAL S6284 : STD_LOGIC;
    SIGNAL S6285 : STD_LOGIC;
    SIGNAL S6286 : STD_LOGIC;
    SIGNAL S6287 : STD_LOGIC;
    SIGNAL S6288 : STD_LOGIC;
    SIGNAL S6289 : STD_LOGIC;
    SIGNAL S6290 : STD_LOGIC;
    SIGNAL S6291 : STD_LOGIC;
    SIGNAL S6292 : STD_LOGIC;
    SIGNAL S6293 : STD_LOGIC;
    SIGNAL S6294 : STD_LOGIC;
    SIGNAL S6295 : STD_LOGIC;
    SIGNAL S6296 : STD_LOGIC;
    SIGNAL S6297 : STD_LOGIC;
    SIGNAL S6298 : STD_LOGIC;
    SIGNAL S6299 : STD_LOGIC;
    SIGNAL S6300 : STD_LOGIC;
    SIGNAL S6301 : STD_LOGIC;
    SIGNAL S6302 : STD_LOGIC;
    SIGNAL S6303 : STD_LOGIC;
    SIGNAL S6304 : STD_LOGIC;
    SIGNAL S6305 : STD_LOGIC;
    SIGNAL S6306 : STD_LOGIC;
    SIGNAL new_controller_1133_S_0 : STD_LOGIC;
    SIGNAL new_controller_1133_Y : STD_LOGIC;
    SIGNAL new_controller_1423_Y_0 : STD_LOGIC;
    SIGNAL new_controller_1423_Y_1 : STD_LOGIC;
    SIGNAL new_controller_234_B_0 : STD_LOGIC;
    SIGNAL new_controller_407_B_0 : STD_LOGIC;
    SIGNAL new_controller_407_B_2 : STD_LOGIC;
    SIGNAL new_controller_clk : STD_LOGIC;
    SIGNAL new_controller_fib_0 : STD_LOGIC;
    SIGNAL new_controller_fib_1 : STD_LOGIC;
    SIGNAL new_controller_fib_2 : STD_LOGIC;
    SIGNAL new_controller_fib_3 : STD_LOGIC;
    SIGNAL new_controller_fib_4 : STD_LOGIC;
    SIGNAL new_controller_opcode_2 : STD_LOGIC;
    SIGNAL new_controller_opcode_3 : STD_LOGIC;
    SIGNAL new_controller_opcode_4 : STD_LOGIC;
    SIGNAL new_controller_opcode_5 : STD_LOGIC;
    SIGNAL new_controller_opcode_6 : STD_LOGIC;
    SIGNAL new_controller_opcode_7 : STD_LOGIC;
    SIGNAL new_controller_outflag_0 : STD_LOGIC;
    SIGNAL new_controller_outflag_1 : STD_LOGIC;
    SIGNAL new_controller_outflag_2 : STD_LOGIC;
    SIGNAL new_controller_outflag_3 : STD_LOGIC;
    SIGNAL new_controller_outflag_6 : STD_LOGIC;
    SIGNAL new_controller_outflag_7 : STD_LOGIC;
    SIGNAL new_controller_pstate_0 : STD_LOGIC;
    SIGNAL new_controller_pstate_1 : STD_LOGIC;
    SIGNAL new_controller_readymem : STD_LOGIC;
    SIGNAL new_controller_rst : STD_LOGIC;
    SIGNAL new_datapath_addrbus_0 : STD_LOGIC;
    SIGNAL new_datapath_addrbus_10 : STD_LOGIC;
    SIGNAL new_datapath_addrbus_11 : STD_LOGIC;
    SIGNAL new_datapath_addrbus_12 : STD_LOGIC;
    SIGNAL new_datapath_addrbus_13 : STD_LOGIC;
    SIGNAL new_datapath_addrbus_14 : STD_LOGIC;
    SIGNAL new_datapath_addrbus_15 : STD_LOGIC;
    SIGNAL new_datapath_addrbus_1 : STD_LOGIC;
    SIGNAL new_datapath_addrbus_2 : STD_LOGIC;
    SIGNAL new_datapath_addrbus_3 : STD_LOGIC;
    SIGNAL new_datapath_addrbus_4 : STD_LOGIC;
    SIGNAL new_datapath_addrbus_5 : STD_LOGIC;
    SIGNAL new_datapath_addrbus_6 : STD_LOGIC;
    SIGNAL new_datapath_addrbus_7 : STD_LOGIC;
    SIGNAL new_datapath_addrbus_8 : STD_LOGIC;
    SIGNAL new_datapath_addrbus_9 : STD_LOGIC;
    SIGNAL new_datapath_addsubunit_in1_0 : STD_LOGIC;
    SIGNAL new_datapath_addsubunit_in1_10 : STD_LOGIC;
    SIGNAL new_datapath_addsubunit_in1_11 : STD_LOGIC;
    SIGNAL new_datapath_addsubunit_in1_12 : STD_LOGIC;
    SIGNAL new_datapath_addsubunit_in1_13 : STD_LOGIC;
    SIGNAL new_datapath_addsubunit_in1_14 : STD_LOGIC;
    SIGNAL new_datapath_addsubunit_in1_15 : STD_LOGIC;
    SIGNAL new_datapath_addsubunit_in1_1 : STD_LOGIC;
    SIGNAL new_datapath_addsubunit_in1_2 : STD_LOGIC;
    SIGNAL new_datapath_addsubunit_in1_3 : STD_LOGIC;
    SIGNAL new_datapath_addsubunit_in1_4 : STD_LOGIC;
    SIGNAL new_datapath_addsubunit_in1_5 : STD_LOGIC;
    SIGNAL new_datapath_addsubunit_in1_6 : STD_LOGIC;
    SIGNAL new_datapath_addsubunit_in1_7 : STD_LOGIC;
    SIGNAL new_datapath_addsubunit_in1_8 : STD_LOGIC;
    SIGNAL new_datapath_addsubunit_in1_9 : STD_LOGIC;
    SIGNAL new_datapath_adr_outreg_0 : STD_LOGIC;
    SIGNAL new_datapath_adr_outreg_10 : STD_LOGIC;
    SIGNAL new_datapath_adr_outreg_11 : STD_LOGIC;
    SIGNAL new_datapath_adr_outreg_12 : STD_LOGIC;
    SIGNAL new_datapath_adr_outreg_13 : STD_LOGIC;
    SIGNAL new_datapath_adr_outreg_14 : STD_LOGIC;
    SIGNAL new_datapath_adr_outreg_15 : STD_LOGIC;
    SIGNAL new_datapath_adr_outreg_1 : STD_LOGIC;
    SIGNAL new_datapath_adr_outreg_2 : STD_LOGIC;
    SIGNAL new_datapath_adr_outreg_3 : STD_LOGIC;
    SIGNAL new_datapath_adr_outreg_4 : STD_LOGIC;
    SIGNAL new_datapath_adr_outreg_5 : STD_LOGIC;
    SIGNAL new_datapath_adr_outreg_6 : STD_LOGIC;
    SIGNAL new_datapath_adr_outreg_7 : STD_LOGIC;
    SIGNAL new_datapath_adr_outreg_8 : STD_LOGIC;
    SIGNAL new_datapath_adr_outreg_9 : STD_LOGIC;
    SIGNAL new_datapath_databusin_0 : STD_LOGIC;
    SIGNAL new_datapath_databusin_10 : STD_LOGIC;
    SIGNAL new_datapath_databusin_11 : STD_LOGIC;
    SIGNAL new_datapath_databusin_12 : STD_LOGIC;
    SIGNAL new_datapath_databusin_13 : STD_LOGIC;
    SIGNAL new_datapath_databusin_14 : STD_LOGIC;
    SIGNAL new_datapath_databusin_15 : STD_LOGIC;
    SIGNAL new_datapath_databusin_1 : STD_LOGIC;
    SIGNAL new_datapath_databusin_2 : STD_LOGIC;
    SIGNAL new_datapath_databusin_3 : STD_LOGIC;
    SIGNAL new_datapath_databusin_4 : STD_LOGIC;
    SIGNAL new_datapath_databusin_5 : STD_LOGIC;
    SIGNAL new_datapath_databusin_6 : STD_LOGIC;
    SIGNAL new_datapath_databusin_7 : STD_LOGIC;
    SIGNAL new_datapath_databusin_8 : STD_LOGIC;
    SIGNAL new_datapath_databusin_9 : STD_LOGIC;
    SIGNAL new_datapath_indatatrf_0 : STD_LOGIC;
    SIGNAL new_datapath_indatatrf_10 : STD_LOGIC;
    SIGNAL new_datapath_indatatrf_11 : STD_LOGIC;
    SIGNAL new_datapath_indatatrf_12 : STD_LOGIC;
    SIGNAL new_datapath_indatatrf_13 : STD_LOGIC;
    SIGNAL new_datapath_indatatrf_14 : STD_LOGIC;
    SIGNAL new_datapath_indatatrf_15 : STD_LOGIC;
    SIGNAL new_datapath_indatatrf_1 : STD_LOGIC;
    SIGNAL new_datapath_indatatrf_2 : STD_LOGIC;
    SIGNAL new_datapath_indatatrf_3 : STD_LOGIC;
    SIGNAL new_datapath_indatatrf_4 : STD_LOGIC;
    SIGNAL new_datapath_indatatrf_5 : STD_LOGIC;
    SIGNAL new_datapath_indatatrf_6 : STD_LOGIC;
    SIGNAL new_datapath_indatatrf_7 : STD_LOGIC;
    SIGNAL new_datapath_indatatrf_8 : STD_LOGIC;
    SIGNAL new_datapath_indatatrf_9 : STD_LOGIC;
    SIGNAL new_datapath_instruction_0 : STD_LOGIC;
    SIGNAL new_datapath_instruction_1 : STD_LOGIC;
    SIGNAL new_datapath_instruction_2 : STD_LOGIC;
    SIGNAL new_datapath_instruction_3 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_1697_B_10 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_1697_B_11 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_1697_B_12 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_1697_B_13 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_1697_B_14 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_1697_B_15 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_1697_B_8 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_1697_B_9 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu1_0 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu1_10 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu1_11 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu1_12 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu1_13 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu1_14 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu1_15 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu1_1 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu1_2 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu1_3 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu1_4 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu1_5 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu1_6 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu1_7 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu1_8 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu1_9 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu2_0 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu2_10 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu2_11 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu2_12 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu2_13 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu2_14 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu2_15 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu2_1 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu2_2 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu2_3 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu2_4 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu2_5 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu2_6 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu2_7 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu2_8 : STD_LOGIC;
    SIGNAL new_datapath_multdivunit_outmdu2_9 : STD_LOGIC;
    SIGNAL new_datapath_muxmem_in2_0 : STD_LOGIC;
    SIGNAL new_datapath_muxmem_in2_10 : STD_LOGIC;
    SIGNAL new_datapath_muxmem_in2_11 : STD_LOGIC;
    SIGNAL new_datapath_muxmem_in2_12 : STD_LOGIC;
    SIGNAL new_datapath_muxmem_in2_13 : STD_LOGIC;
    SIGNAL new_datapath_muxmem_in2_14 : STD_LOGIC;
    SIGNAL new_datapath_muxmem_in2_15 : STD_LOGIC;
    SIGNAL new_datapath_muxmem_in2_1 : STD_LOGIC;
    SIGNAL new_datapath_muxmem_in2_2 : STD_LOGIC;
    SIGNAL new_datapath_muxmem_in2_3 : STD_LOGIC;
    SIGNAL new_datapath_muxmem_in2_4 : STD_LOGIC;
    SIGNAL new_datapath_muxmem_in2_5 : STD_LOGIC;
    SIGNAL new_datapath_muxmem_in2_6 : STD_LOGIC;
    SIGNAL new_datapath_muxmem_in2_7 : STD_LOGIC;
    SIGNAL new_datapath_muxmem_in2_8 : STD_LOGIC;
    SIGNAL new_datapath_muxmem_in2_9 : STD_LOGIC;
    SIGNAL new_datapath_muxrd_outmux_0 : STD_LOGIC;
    SIGNAL new_datapath_muxrd_outmux_1 : STD_LOGIC;
    SIGNAL new_datapath_muxrd_outmux_2 : STD_LOGIC;
    SIGNAL new_datapath_muxrd_outmux_3 : STD_LOGIC;
    SIGNAL new_datapath_muxrs1_outmux_0 : STD_LOGIC;
    SIGNAL new_datapath_muxrs1_outmux_1 : STD_LOGIC;
    SIGNAL new_datapath_muxrs1_outmux_2 : STD_LOGIC;
    SIGNAL new_datapath_muxrs1_outmux_3 : STD_LOGIC;
    SIGNAL new_datapath_muxrs2_outmux_0 : STD_LOGIC;
    SIGNAL new_datapath_muxrs2_outmux_1 : STD_LOGIC;
    SIGNAL new_datapath_muxrs2_outmux_2 : STD_LOGIC;
    SIGNAL new_datapath_muxrs2_outmux_3 : STD_LOGIC;
    SIGNAL new_datapath_p1trf_0 : STD_LOGIC;
    SIGNAL new_datapath_p1trf_1 : STD_LOGIC;
    SIGNAL new_datapath_p1trf_2 : STD_LOGIC;
    SIGNAL new_datapath_p1trf_3 : STD_LOGIC;
    SIGNAL new_datapath_p1trf_4 : STD_LOGIC;
    SIGNAL new_datapath_p1trf_5 : STD_LOGIC;
    SIGNAL new_datapath_p1trf_6 : STD_LOGIC;
    SIGNAL new_datapath_p1trf_7 : STD_LOGIC;
    SIGNAL new_datapath_p2trf_0 : STD_LOGIC;
    SIGNAL new_datapath_p2trf_1 : STD_LOGIC;
    SIGNAL new_datapath_p2trf_2 : STD_LOGIC;
    SIGNAL new_datapath_p2trf_3 : STD_LOGIC;
    SIGNAL new_datapath_p2trf_4 : STD_LOGIC;
    SIGNAL new_datapath_p2trf_5 : STD_LOGIC;
    SIGNAL new_datapath_p2trf_6 : STD_LOGIC;
    SIGNAL new_datapath_p2trf_7 : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_1961_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_1979_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_1997_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2015_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2033_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2051_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2069_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2087_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2105_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2123_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2141_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2159_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2177_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2195_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2213_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2231_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2265_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2283_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2301_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2319_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2337_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2355_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2373_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2391_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2409_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2427_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2445_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2463_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2481_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2499_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2517_A : STD_LOGIC;
    SIGNAL new_datapath_shiftunit_2534_A : STD_LOGIC;

BEGIN
notg_0: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_outmdu2_15,
        out1 => S2581
    );
notg_1: ENTITY WORK.notg
    PORT MAP (
        in1 => new_controller_opcode_7,
        out1 => S2592
    );
notg_2: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_databusin_15,
        out1 => S2603
    );
notg_3: ENTITY WORK.notg
    PORT MAP (
        in1 => new_controller_outflag_7,
        out1 => S2614
    );
notg_4: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_muxmem_in2_0,
        out1 => S2625
    );
notg_5: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_muxmem_in2_1,
        out1 => S2636
    );
notg_6: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_muxmem_in2_2,
        out1 => S2647
    );
notg_7: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_muxmem_in2_3,
        out1 => S2658
    );
notg_8: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_muxmem_in2_4,
        out1 => S2669
    );
notg_9: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_muxmem_in2_5,
        out1 => S2680
    );
notg_10: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_muxmem_in2_6,
        out1 => S2690
    );
notg_11: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_muxmem_in2_7,
        out1 => S2701
    );
notg_12: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_muxmem_in2_8,
        out1 => S2712
    );
notg_13: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_muxmem_in2_9,
        out1 => S2723
    );
notg_14: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_muxmem_in2_10,
        out1 => S2734
    );
notg_15: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_muxmem_in2_11,
        out1 => S2745
    );
notg_16: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_muxmem_in2_12,
        out1 => S2756
    );
notg_17: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_muxmem_in2_13,
        out1 => S2767
    );
notg_18: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_muxmem_in2_14,
        out1 => S2778
    );
notg_19: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_outmdu1_6,
        out1 => S2789
    );
notg_20: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_outmdu2_0,
        out1 => S2800
    );
notg_21: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_outmdu2_1,
        out1 => S2811
    );
notg_22: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_outmdu2_2,
        out1 => S2822
    );
notg_23: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_outmdu2_3,
        out1 => S2832
    );
notg_24: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_outmdu2_4,
        out1 => S2843
    );
notg_25: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_outmdu2_5,
        out1 => S2854
    );
notg_26: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_outmdu2_6,
        out1 => S2865
    );
notg_27: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_outmdu2_7,
        out1 => S2876
    );
notg_28: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_outmdu2_8,
        out1 => S2887
    );
notg_29: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_outmdu2_9,
        out1 => S2898
    );
notg_30: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_outmdu2_10,
        out1 => S2909
    );
notg_31: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_outmdu2_11,
        out1 => S2920
    );
notg_32: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_outmdu2_12,
        out1 => S2931
    );
notg_33: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_outmdu2_13,
        out1 => S2942
    );
notg_34: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_outmdu2_14,
        out1 => S2953
    );
notg_35: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_instruction_0,
        out1 => S2964
    );
notg_36: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_instruction_3,
        out1 => S2975
    );
notg_37: ENTITY WORK.notg
    PORT MAP (
        in1 => new_controller_fib_0,
        out1 => S2985
    );
notg_38: ENTITY WORK.notg
    PORT MAP (
        in1 => new_controller_fib_1,
        out1 => S2996
    );
notg_39: ENTITY WORK.notg
    PORT MAP (
        in1 => new_controller_fib_2,
        out1 => S3007
    );
notg_40: ENTITY WORK.notg
    PORT MAP (
        in1 => new_controller_fib_3,
        out1 => S3018
    );
notg_41: ENTITY WORK.notg
    PORT MAP (
        in1 => new_controller_fib_4,
        out1 => S3029
    );
notg_42: ENTITY WORK.notg
    PORT MAP (
        in1 => new_controller_234_B_0,
        out1 => S3040
    );
notg_43: ENTITY WORK.notg
    PORT MAP (
        in1 => new_controller_opcode_2,
        out1 => S3051
    );
notg_44: ENTITY WORK.notg
    PORT MAP (
        in1 => new_controller_opcode_3,
        out1 => S3062
    );
notg_45: ENTITY WORK.notg
    PORT MAP (
        in1 => new_controller_opcode_4,
        out1 => S3073
    );
notg_46: ENTITY WORK.notg
    PORT MAP (
        in1 => new_controller_opcode_5,
        out1 => S3084
    );
notg_47: ENTITY WORK.notg
    PORT MAP (
        in1 => new_controller_opcode_6,
        out1 => S3095
    );
notg_48: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_databusin_14,
        out1 => S3106
    );
notg_49: ENTITY WORK.notg
    PORT MAP (
        in1 => new_controller_407_B_0,
        out1 => S3117
    );
notg_50: ENTITY WORK.notg
    PORT MAP (
        in1 => new_controller_pstate_1,
        out1 => S3128
    );
notg_51: ENTITY WORK.notg
    PORT MAP (
        in1 => new_controller_pstate_0,
        out1 => S3139
    );
notg_52: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_p1trf_0,
        out1 => S3150
    );
notg_53: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_p1trf_1,
        out1 => S3160
    );
notg_54: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_p1trf_2,
        out1 => S3171
    );
notg_55: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_p1trf_3,
        out1 => S3182
    );
notg_56: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_p1trf_4,
        out1 => S3193
    );
notg_57: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_p1trf_5,
        out1 => S3204
    );
notg_58: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_p1trf_6,
        out1 => S3215
    );
notg_59: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_p1trf_7,
        out1 => S3226
    );
notg_60: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_p2trf_0,
        out1 => S3237
    );
notg_61: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_p2trf_1,
        out1 => S3248
    );
notg_62: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_p2trf_2,
        out1 => S3259
    );
notg_63: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_p2trf_3,
        out1 => S3270
    );
notg_64: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_p2trf_4,
        out1 => S3281
    );
notg_65: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_p2trf_5,
        out1 => S3292
    );
notg_66: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_p2trf_6,
        out1 => S3303
    );
notg_67: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_p2trf_7,
        out1 => S3314
    );
notg_68: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_8,
        out1 => S3325
    );
notg_69: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_9,
        out1 => S3336
    );
notg_70: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_10,
        out1 => S3346
    );
notg_71: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_11,
        out1 => S3357
    );
notg_72: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_12,
        out1 => S3368
    );
notg_73: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_13,
        out1 => S3379
    );
notg_74: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_14,
        out1 => S3390
    );
notg_75: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_15,
        out1 => S3401
    );
notg_76: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_1697_B_14,
        out1 => S3412
    );
notg_77: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_1697_B_13,
        out1 => S3423
    );
notg_78: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_1697_B_12,
        out1 => S3434
    );
notg_79: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_1697_B_11,
        out1 => S3445
    );
notg_80: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_1697_B_10,
        out1 => S3456
    );
notg_81: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_1697_B_9,
        out1 => S3467
    );
notg_82: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_multdivunit_1697_B_8,
        out1 => S3478
    );
notg_83: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_shiftunit_1997_A,
        out1 => S3489
    );
notg_84: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_shiftunit_2015_A,
        out1 => S3500
    );
notg_85: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_shiftunit_2069_A,
        out1 => S3511
    );
notg_86: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_shiftunit_2087_A,
        out1 => S3522
    );
notg_87: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_shiftunit_2105_A,
        out1 => S3533
    );
notg_88: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_shiftunit_2123_A,
        out1 => S3544
    );
notg_89: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_shiftunit_2141_A,
        out1 => S3554
    );
notg_90: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_shiftunit_2159_A,
        out1 => S3565
    );
notg_91: ENTITY WORK.notg
    PORT MAP (
        in1 => new_datapath_shiftunit_2177_A,
        out1 => S3576
    );
nor_n_92: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_controller_opcode_6,
        in1(1) => new_controller_opcode_7,
        out1 => S3587
    );
notg_93: ENTITY WORK.notg
    PORT MAP (
        in1 => S3587,
        out1 => S3598
    );
nor_n_94: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3084,
        in1(1) => new_controller_opcode_4,
        out1 => S3609
    );
nand_n_95: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_opcode_5,
        in1(1) => S3073,
        out1 => S3620
    );
nor_n_96: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3598,
        in1(1) => new_controller_opcode_4,
        out1 => S3631
    );
nor_n_97: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3620,
        in1(1) => S3598,
        out1 => S3642
    );
nand_n_98: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3609,
        in1(1) => S3587,
        out1 => S3653
    );
nor_n_99: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_controller_pstate_0,
        in1(1) => S3128,
        out1 => S3664
    );
notg_100: ENTITY WORK.notg
    PORT MAP (
        in1 => S3664,
        out1 => S3675
    );
nor_n_101: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3653,
        in1(1) => new_controller_opcode_3,
        out1 => S3686
    );
notg_102: ENTITY WORK.notg
    PORT MAP (
        in1 => S3686,
        out1 => S3697
    );
nor_n_103: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3697,
        in1(1) => S3675,
        out1 => S3708
    );
nand_n_104: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3686,
        in1(1) => S3664,
        out1 => S3719
    );
nor_n_105: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3719,
        in1(1) => new_controller_opcode_2,
        out1 => S6215
    );
notg_106: ENTITY WORK.notg
    PORT MAP (
        in1 => S6215,
        out1 => S3740
    );
nor_n_107: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3719,
        in1(1) => S3051,
        out1 => S6216
    );
nor_n_108: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3139,
        in1(1) => new_controller_pstate_1,
        out1 => S3761
    );
nand_n_109: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_pstate_0,
        in1(1) => S3128,
        out1 => S3771
    );
nand_n_110: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_opcode_6,
        in1(1) => new_controller_opcode_7,
        out1 => S3782
    );
notg_111: ENTITY WORK.notg
    PORT MAP (
        in1 => S3782,
        out1 => S3793
    );
nor_n_112: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3793,
        in1(1) => S3631,
        out1 => S3804
    );
nor_n_113: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3084,
        in1(1) => S3073,
        out1 => S3815
    );
nand_n_114: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_opcode_5,
        in1(1) => new_controller_opcode_4,
        out1 => S3826
    );
nor_n_115: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3826,
        in1(1) => S3782,
        out1 => S3837
    );
nor_n_116: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3062,
        in1(1) => new_controller_opcode_2,
        out1 => S3848
    );
nand_n_117: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_opcode_3,
        in1(1) => S3051,
        out1 => S3859
    );
nand_n_118: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3837,
        in1(1) => new_controller_opcode_3,
        out1 => S3870
    );
nor_n_119: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3870,
        in1(1) => new_controller_opcode_2,
        out1 => S3881
    );
notg_120: ENTITY WORK.notg
    PORT MAP (
        in1 => S3881,
        out1 => S3892
    );
nor_n_121: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_controller_opcode_5,
        in1(1) => new_controller_opcode_4,
        out1 => S3903
    );
nand_n_122: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3084,
        in1(1) => S3073,
        out1 => S3914
    );
nor_n_123: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3903,
        in1(1) => S3804,
        out1 => S3925
    );
nand_n_124: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3925,
        in1(1) => S3892,
        out1 => S3936
    );
nand_n_125: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3642,
        in1(1) => new_controller_opcode_3,
        out1 => S3947
    );
nand_n_126: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3859,
        in1(1) => S3837,
        out1 => S3958
    );
nor_n_127: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_controller_opcode_3,
        in1(1) => S3051,
        out1 => S3969
    );
nand_n_128: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3969,
        in1(1) => new_controller_fib_2,
        out1 => S3980
    );
nor_n_129: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3980,
        in1(1) => S2996,
        out1 => S3990
    );
nor_n_130: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3990,
        in1(1) => S3958,
        out1 => S4001
    );
notg_131: ENTITY WORK.notg
    PORT MAP (
        in1 => S4001,
        out1 => S4012
    );
nand_n_132: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4012,
        in1(1) => S3947,
        out1 => S4023
    );
nor_n_133: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4023,
        in1(1) => S3936,
        out1 => S4034
    );
nor_n_134: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4034,
        in1(1) => S3771,
        out1 => S4045
    );
nor_n_135: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_controller_opcode_5,
        in1(1) => S3073,
        out1 => S4056
    );
nand_n_136: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3084,
        in1(1) => new_controller_opcode_4,
        out1 => S4067
    );
nor_n_137: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4056,
        in1(1) => S3609,
        out1 => S4078
    );
nand_n_138: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4067,
        in1(1) => S3620,
        out1 => S4089
    );
nor_n_139: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4078,
        in1(1) => S3782,
        out1 => S4100
    );
notg_140: ENTITY WORK.notg
    PORT MAP (
        in1 => S4100,
        out1 => S4111
    );
nor_n_141: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4111,
        in1(1) => S3128,
        out1 => S4122
    );
nand_n_142: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4100,
        in1(1) => new_controller_pstate_1,
        out1 => S4133
    );
nor_n_143: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4133,
        in1(1) => S3139,
        out1 => S4144
    );
nand_n_144: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4122,
        in1(1) => new_controller_pstate_0,
        out1 => S4155
    );
nor_n_145: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_controller_readymem,
        in1(1) => new_controller_234_B_0,
        out1 => S4166
    );
notg_146: ENTITY WORK.notg
    PORT MAP (
        in1 => S4166,
        out1 => S4177
    );
nand_n_147: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4177,
        in1(1) => S3708,
        out1 => S4188
    );
nand_n_148: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4188,
        in1(1) => S4155,
        out1 => S4199
    );
nor_n_149: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4199,
        in1(1) => S4045,
        out1 => S4210
    );
nand_n_150: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4210,
        in1(1) => new_datapath_muxmem_in2_15,
        out1 => S4221
    );
nand_n_151: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3761,
        in1(1) => S3609,
        out1 => S4232
    );
notg_152: ENTITY WORK.notg
    PORT MAP (
        in1 => S4232,
        out1 => S4237
    );
nor_n_153: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3771,
        in1(1) => S3653,
        out1 => S4238
    );
nand_n_154: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3761,
        in1(1) => S3642,
        out1 => S4246
    );
nor_n_155: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4246,
        in1(1) => S3062,
        out1 => S4254
    );
nand_n_156: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4238,
        in1(1) => new_controller_opcode_3,
        out1 => S4261
    );
nand_n_157: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_opcode_3,
        in1(1) => new_controller_opcode_2,
        out1 => S4269
    );
notg_158: ENTITY WORK.notg
    PORT MAP (
        in1 => S4269,
        out1 => S4278
    );
nor_n_159: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4269,
        in1(1) => S4246,
        out1 => S4289
    );
nand_n_160: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4289,
        in1(1) => new_controller_234_B_0,
        out1 => S4300
    );
nand_n_161: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4269,
        in1(1) => S4238,
        out1 => S4311
    );
nor_n_162: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_controller_407_B_2,
        in1(1) => new_controller_fib_0,
        out1 => S4322
    );
notg_163: ENTITY WORK.notg
    PORT MAP (
        in1 => S4322,
        out1 => S4333
    );
nor_n_164: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_controller_407_B_2,
        in1(1) => new_controller_407_B_0,
        out1 => S4344
    );
nor_n_165: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_controller_fib_2,
        in1(1) => S2996,
        out1 => S4355
    );
nand_n_166: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4355,
        in1(1) => S4333,
        out1 => S4366
    );
nor_n_167: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4366,
        in1(1) => S4344,
        out1 => S4377
    );
nor_n_168: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_controller_fib_1,
        in1(1) => new_controller_fib_0,
        out1 => S4388
    );
nand_n_169: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4388,
        in1(1) => new_controller_fib_2,
        out1 => S4399
    );
notg_170: ENTITY WORK.notg
    PORT MAP (
        in1 => S4399,
        out1 => S4410
    );
nor_n_171: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_controller_fib_2,
        in1(1) => S2985,
        out1 => S4421
    );
nand_n_172: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3007,
        in1(1) => new_controller_fib_0,
        out1 => S4432
    );
nor_n_173: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4432,
        in1(1) => new_controller_fib_1,
        out1 => S4443
    );
nor_n_174: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4443,
        in1(1) => S4410,
        out1 => S4454
    );
nor_n_175: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4454,
        in1(1) => new_controller_407_B_2,
        out1 => S4465
    );
nor_n_176: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4465,
        in1(1) => new_controller_407_B_0,
        out1 => S4476
    );
nand_n_177: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4388,
        in1(1) => S3007,
        out1 => S4487
    );
nor_n_178: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4388,
        in1(1) => S3117,
        out1 => S4498
    );
nor_n_179: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4498,
        in1(1) => S4476,
        out1 => S4509
    );
nor_n_180: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4509,
        in1(1) => S4377,
        out1 => S4519
    );
notg_181: ENTITY WORK.notg
    PORT MAP (
        in1 => S4519,
        out1 => S4530
    );
nand_n_182: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3969,
        in1(1) => new_controller_234_B_0,
        out1 => S4541
    );
nor_n_183: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3782,
        in1(1) => S3771,
        out1 => S4552
    );
nand_n_184: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3793,
        in1(1) => S3761,
        out1 => S4563
    );
nor_n_185: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4563,
        in1(1) => S3826,
        out1 => S4570
    );
nand_n_186: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3837,
        in1(1) => S3761,
        out1 => S4578
    );
nor_n_187: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4578,
        in1(1) => S4541,
        out1 => S4586
    );
nand_n_188: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4586,
        in1(1) => S4530,
        out1 => S4593
    );
nand_n_189: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4593,
        in1(1) => S4311,
        out1 => S4602
    );
nand_n_190: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4602,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S4613
    );
nand_n_191: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4613,
        in1(1) => S4300,
        out1 => S4621
    );
nand_n_192: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4621,
        in1(1) => new_datapath_muxmem_in2_14,
        out1 => S4632
    );
notg_193: ENTITY WORK.notg
    PORT MAP (
        in1 => S4632,
        out1 => S4643
    );
nor_n_194: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4621,
        in1(1) => new_datapath_muxmem_in2_14,
        out1 => S4654
    );
nor_n_195: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4654,
        in1(1) => S4643,
        out1 => S4665
    );
nand_n_196: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4602,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S4676
    );
nand_n_197: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4676,
        in1(1) => S4300,
        out1 => S4686
    );
nand_n_198: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4686,
        in1(1) => new_datapath_muxmem_in2_13,
        out1 => S4697
    );
notg_199: ENTITY WORK.notg
    PORT MAP (
        in1 => S4697,
        out1 => S4708
    );
nor_n_200: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4686,
        in1(1) => new_datapath_muxmem_in2_13,
        out1 => S4718
    );
nand_n_201: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4602,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S4729
    );
nand_n_202: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4729,
        in1(1) => S4300,
        out1 => S4740
    );
nand_n_203: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4740,
        in1(1) => new_datapath_muxmem_in2_12,
        out1 => S4750
    );
notg_204: ENTITY WORK.notg
    PORT MAP (
        in1 => S4750,
        out1 => S4761
    );
nor_n_205: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4740,
        in1(1) => new_datapath_muxmem_in2_12,
        out1 => S4772
    );
nor_n_206: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4772,
        in1(1) => S4761,
        out1 => S4783
    );
nand_n_207: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4602,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S4793
    );
nand_n_208: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4793,
        in1(1) => S4300,
        out1 => S4804
    );
notg_209: ENTITY WORK.notg
    PORT MAP (
        in1 => S4804,
        out1 => S4815
    );
nor_n_210: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4804,
        in1(1) => new_datapath_muxmem_in2_11,
        out1 => S4825
    );
nor_n_211: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4815,
        in1(1) => S2745,
        out1 => S4836
    );
nand_n_212: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4602,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S4847
    );
nand_n_213: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4847,
        in1(1) => S4300,
        out1 => S4857
    );
nand_n_214: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4857,
        in1(1) => new_datapath_muxmem_in2_10,
        out1 => S4868
    );
notg_215: ENTITY WORK.notg
    PORT MAP (
        in1 => S4868,
        out1 => S4879
    );
nor_n_216: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4857,
        in1(1) => new_datapath_muxmem_in2_10,
        out1 => S4890
    );
nor_n_217: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4890,
        in1(1) => S4879,
        out1 => S4900
    );
nand_n_218: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4602,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S4911
    );
nand_n_219: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4911,
        in1(1) => S4300,
        out1 => S4922
    );
nand_n_220: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4922,
        in1(1) => new_datapath_muxmem_in2_9,
        out1 => S4932
    );
notg_221: ENTITY WORK.notg
    PORT MAP (
        in1 => S4932,
        out1 => S4943
    );
nor_n_222: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4922,
        in1(1) => new_datapath_muxmem_in2_9,
        out1 => S4954
    );
nand_n_223: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4602,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S4964
    );
nand_n_224: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4964,
        in1(1) => S4300,
        out1 => S4975
    );
nand_n_225: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4975,
        in1(1) => new_datapath_muxmem_in2_8,
        out1 => S4986
    );
notg_226: ENTITY WORK.notg
    PORT MAP (
        in1 => S4986,
        out1 => S4997
    );
nor_n_227: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4975,
        in1(1) => new_datapath_muxmem_in2_8,
        out1 => S5007
    );
nor_n_228: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5007,
        in1(1) => S4997,
        out1 => S5018
    );
nor_n_229: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_controller_fib_1,
        in1(1) => S2985,
        out1 => S5029
    );
nand_n_230: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_fib_2,
        in1(1) => new_controller_fib_0,
        out1 => S5039
    );
nor_n_231: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5039,
        in1(1) => new_controller_fib_1,
        out1 => S5050
    );
nand_n_232: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5029,
        in1(1) => new_controller_fib_2,
        out1 => S5061
    );
nand_n_233: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5050,
        in1(1) => S3117,
        out1 => S5072
    );
nand_n_234: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5072,
        in1(1) => S4519,
        out1 => S5082
    );
notg_235: ENTITY WORK.notg
    PORT MAP (
        in1 => S5082,
        out1 => S5093
    );
nand_n_236: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4238,
        in1(1) => S3969,
        out1 => S5104
    );
nor_n_237: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3892,
        in1(1) => S3771,
        out1 => S5115
    );
nand_n_238: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3881,
        in1(1) => S3761,
        out1 => S5125
    );
nor_n_239: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3095,
        in1(1) => new_controller_opcode_7,
        out1 => S5136
    );
nand_n_240: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_opcode_6,
        in1(1) => S2592,
        out1 => S5147
    );
nor_n_241: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5147,
        in1(1) => S4232,
        out1 => S5157
    );
nand_n_242: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5136,
        in1(1) => S4237,
        out1 => S5168
    );
nor_n_243: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5157,
        in1(1) => S5115,
        out1 => S5179
    );
nand_n_244: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5179,
        in1(1) => S5104,
        out1 => S5190
    );
nor_n_245: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3969,
        in1(1) => S3848,
        out1 => S5200
    );
nand_n_246: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5200,
        in1(1) => S4570,
        out1 => S5211
    );
notg_247: ENTITY WORK.notg
    PORT MAP (
        in1 => S5211,
        out1 => S5222
    );
nand_n_248: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5222,
        in1(1) => new_controller_234_B_0,
        out1 => S5232
    );
nor_n_249: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5147,
        in1(1) => S3914,
        out1 => S5239
    );
nand_n_250: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5136,
        in1(1) => S3903,
        out1 => S5247
    );
nor_n_251: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3914,
        in1(1) => S3782,
        out1 => S5255
    );
nand_n_252: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3903,
        in1(1) => S3793,
        out1 => S5262
    );
nor_n_253: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_controller_opcode_6,
        in1(1) => S2592,
        out1 => S5271
    );
nand_n_254: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3095,
        in1(1) => new_controller_opcode_7,
        out1 => S5280
    );
nor_n_255: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5280,
        in1(1) => S3826,
        out1 => S5290
    );
nand_n_256: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5271,
        in1(1) => S3815,
        out1 => S5300
    );
nor_n_257: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5290,
        in1(1) => S5255,
        out1 => S5311
    );
nand_n_258: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5300,
        in1(1) => S5262,
        out1 => S5322
    );
nand_n_259: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5311,
        in1(1) => S5247,
        out1 => S5332
    );
nand_n_260: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5322,
        in1(1) => S3761,
        out1 => S5343
    );
nand_n_261: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5332,
        in1(1) => S3761,
        out1 => S5354
    );
notg_262: ENTITY WORK.notg
    PORT MAP (
        in1 => S5354,
        out1 => S5365
    );
nand_n_263: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5354,
        in1(1) => S5232,
        out1 => S5376
    );
nor_n_264: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5376,
        in1(1) => S5190,
        out1 => S5387
    );
nor_n_265: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5093,
        in1(1) => S4578,
        out1 => S5398
    );
nand_n_266: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5398,
        in1(1) => S3969,
        out1 => S5408
    );
notg_267: ENTITY WORK.notg
    PORT MAP (
        in1 => S5408,
        out1 => S5419
    );
nand_n_268: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5408,
        in1(1) => S5387,
        out1 => S5430
    );
nand_n_269: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5430,
        in1(1) => new_datapath_instruction_3,
        out1 => S5440
    );
nor_n_270: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3826,
        in1(1) => S3598,
        out1 => S5451
    );
nand_n_271: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3815,
        in1(1) => S3587,
        out1 => S5462
    );
nor_n_272: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5280,
        in1(1) => S4078,
        out1 => S5473
    );
nand_n_273: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5271,
        in1(1) => S4089,
        out1 => S5483
    );
nor_n_274: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5473,
        in1(1) => S5451,
        out1 => S5494
    );
nand_n_275: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5483,
        in1(1) => S5462,
        out1 => S5505
    );
nor_n_276: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5494,
        in1(1) => S3771,
        out1 => S5515
    );
nand_n_277: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5505,
        in1(1) => S3761,
        out1 => S5526
    );
nor_n_278: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4563,
        in1(1) => S3620,
        out1 => S5537
    );
nand_n_279: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4552,
        in1(1) => S3609,
        out1 => S5547
    );
nand_n_280: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3761,
        in1(1) => new_controller_opcode_4,
        out1 => S5558
    );
notg_281: ENTITY WORK.notg
    PORT MAP (
        in1 => S5558,
        out1 => S5568
    );
nor_n_282: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4563,
        in1(1) => S4067,
        out1 => S5579
    );
nand_n_283: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4552,
        in1(1) => S4056,
        out1 => S5590
    );
nor_n_284: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4563,
        in1(1) => S4078,
        out1 => S5600
    );
nand_n_285: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4552,
        in1(1) => S4089,
        out1 => S5611
    );
nor_n_286: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5280,
        in1(1) => S3914,
        out1 => S5621
    );
nand_n_287: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5271,
        in1(1) => S3903,
        out1 => S5632
    );
nor_n_288: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5147,
        in1(1) => S3826,
        out1 => S5642
    );
nand_n_289: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5136,
        in1(1) => S3815,
        out1 => S5653
    );
nor_n_290: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5642,
        in1(1) => S5621,
        out1 => S5663
    );
nand_n_291: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5653,
        in1(1) => S5632,
        out1 => S5673
    );
nor_n_292: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5663,
        in1(1) => S3771,
        out1 => S5683
    );
nand_n_293: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5673,
        in1(1) => S3761,
        out1 => S5693
    );
nor_n_294: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5683,
        in1(1) => S5600,
        out1 => S5702
    );
nand_n_295: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5693,
        in1(1) => S5611,
        out1 => S5710
    );
nor_n_296: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5710,
        in1(1) => S5515,
        out1 => S5719
    );
nand_n_297: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5702,
        in1(1) => S5526,
        out1 => S5729
    );
nor_n_298: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4246,
        in1(1) => new_controller_opcode_2,
        out1 => S5739
    );
nor_n_299: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5739,
        in1(1) => S6216,
        out1 => S5749
    );
nor_n_300: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5211,
        in1(1) => new_controller_234_B_0,
        out1 => S5759
    );
nor_n_301: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5759,
        in1(1) => S5729,
        out1 => S5770
    );
nand_n_302: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5770,
        in1(1) => S5749,
        out1 => S5780
    );
nand_n_303: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5780,
        in1(1) => new_controller_fib_3,
        out1 => S5791
    );
nand_n_304: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5791,
        in1(1) => S5440,
        out1 => new_datapath_muxrs1_outmux_3
    );
nand_n_305: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5430,
        in1(1) => new_datapath_instruction_0,
        out1 => S5810
    );
nand_n_306: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5780,
        in1(1) => new_controller_fib_0,
        out1 => S5821
    );
nand_n_307: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5821,
        in1(1) => S5810,
        out1 => new_datapath_muxrs1_outmux_0
    );
nand_n_308: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_muxrs1_outmux_0,
        in1(1) => new_datapath_muxrs1_outmux_3,
        out1 => S5841
    );
nand_n_309: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5430,
        in1(1) => new_datapath_instruction_1,
        out1 => S5852
    );
nand_n_310: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5780,
        in1(1) => new_controller_fib_1,
        out1 => S5862
    );
nand_n_311: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5862,
        in1(1) => S5852,
        out1 => new_datapath_muxrs1_outmux_1
    );
nand_n_312: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5430,
        in1(1) => new_datapath_instruction_2,
        out1 => S5882
    );
nand_n_313: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5780,
        in1(1) => new_controller_fib_2,
        out1 => S5893
    );
nand_n_314: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5893,
        in1(1) => S5882,
        out1 => new_datapath_muxrs1_outmux_2
    );
nand_n_315: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_muxrs1_outmux_2,
        in1(1) => new_datapath_muxrs1_outmux_1,
        out1 => S5902
    );
nor_n_316: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5902,
        in1(1) => S5841,
        out1 => S5903
    );
nand_n_317: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5903,
        in1(1) => new_controller_outflag_7,
        out1 => S5904
    );
notg_318: ENTITY WORK.notg
    PORT MAP (
        in1 => S5904,
        out1 => S5905
    );
nor_n_319: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5903,
        in1(1) => S3226,
        out1 => S5906
    );
nor_n_320: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5906,
        in1(1) => S5905,
        out1 => S5907
    );
notg_321: ENTITY WORK.notg
    PORT MAP (
        in1 => S5907,
        out1 => new_datapath_addsubunit_in1_7
    );
nand_n_322: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_7,
        in1(1) => S4602,
        out1 => S5908
    );
nand_n_323: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5908,
        in1(1) => S4300,
        out1 => S5909
    );
nand_n_324: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5909,
        in1(1) => new_datapath_muxmem_in2_7,
        out1 => S5910
    );
notg_325: ENTITY WORK.notg
    PORT MAP (
        in1 => S5910,
        out1 => S5911
    );
nor_n_326: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5909,
        in1(1) => new_datapath_muxmem_in2_7,
        out1 => S5912
    );
nand_n_327: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5903,
        in1(1) => new_controller_outflag_6,
        out1 => S5913
    );
notg_328: ENTITY WORK.notg
    PORT MAP (
        in1 => S5913,
        out1 => S5914
    );
nor_n_329: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5903,
        in1(1) => S3215,
        out1 => S5915
    );
nor_n_330: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5915,
        in1(1) => S5914,
        out1 => S5916
    );
notg_331: ENTITY WORK.notg
    PORT MAP (
        in1 => S5916,
        out1 => new_datapath_addsubunit_in1_6
    );
nand_n_332: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_6,
        in1(1) => S4602,
        out1 => S5917
    );
nand_n_333: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5917,
        in1(1) => S4300,
        out1 => S5918
    );
nand_n_334: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5918,
        in1(1) => new_datapath_muxmem_in2_6,
        out1 => S5919
    );
notg_335: ENTITY WORK.notg
    PORT MAP (
        in1 => S5919,
        out1 => S5920
    );
nor_n_336: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5918,
        in1(1) => new_datapath_muxmem_in2_6,
        out1 => S5921
    );
nor_n_337: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5921,
        in1(1) => S5920,
        out1 => S5922
    );
nand_n_338: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5903,
        in1(1) => new_controller_407_B_2,
        out1 => S5923
    );
notg_339: ENTITY WORK.notg
    PORT MAP (
        in1 => S5923,
        out1 => S5924
    );
nor_n_340: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5903,
        in1(1) => S3204,
        out1 => S5925
    );
nor_n_341: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5925,
        in1(1) => S5924,
        out1 => S5926
    );
notg_342: ENTITY WORK.notg
    PORT MAP (
        in1 => S5926,
        out1 => new_datapath_addsubunit_in1_5
    );
nand_n_343: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_5,
        in1(1) => S4602,
        out1 => S5927
    );
nand_n_344: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5927,
        in1(1) => S4300,
        out1 => S5928
    );
nand_n_345: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5928,
        in1(1) => new_datapath_muxmem_in2_5,
        out1 => S5929
    );
notg_346: ENTITY WORK.notg
    PORT MAP (
        in1 => S5929,
        out1 => S5930
    );
nor_n_347: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5928,
        in1(1) => new_datapath_muxmem_in2_5,
        out1 => S5931
    );
nand_n_348: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4289,
        in1(1) => new_controller_fib_4,
        out1 => S5932
    );
nand_n_349: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5903,
        in1(1) => new_controller_407_B_0,
        out1 => S5933
    );
notg_350: ENTITY WORK.notg
    PORT MAP (
        in1 => S5933,
        out1 => S5934
    );
nor_n_351: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5903,
        in1(1) => S3193,
        out1 => S5935
    );
nor_n_352: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5935,
        in1(1) => S5934,
        out1 => S5936
    );
notg_353: ENTITY WORK.notg
    PORT MAP (
        in1 => S5936,
        out1 => new_datapath_addsubunit_in1_4
    );
nand_n_354: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_4,
        in1(1) => S4602,
        out1 => S5937
    );
nand_n_355: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5937,
        in1(1) => S5932,
        out1 => S5938
    );
nand_n_356: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5938,
        in1(1) => new_datapath_muxmem_in2_4,
        out1 => S5939
    );
notg_357: ENTITY WORK.notg
    PORT MAP (
        in1 => S5939,
        out1 => S5940
    );
nor_n_358: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5938,
        in1(1) => new_datapath_muxmem_in2_4,
        out1 => S5941
    );
nor_n_359: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5941,
        in1(1) => S5940,
        out1 => S5942
    );
nand_n_360: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4289,
        in1(1) => new_controller_fib_3,
        out1 => S5943
    );
nand_n_361: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5903,
        in1(1) => new_controller_outflag_3,
        out1 => S5944
    );
notg_362: ENTITY WORK.notg
    PORT MAP (
        in1 => S5944,
        out1 => S5945
    );
nor_n_363: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5903,
        in1(1) => S3182,
        out1 => S5946
    );
nor_n_364: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5946,
        in1(1) => S5945,
        out1 => S5947
    );
notg_365: ENTITY WORK.notg
    PORT MAP (
        in1 => S5947,
        out1 => new_datapath_addsubunit_in1_3
    );
nand_n_366: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_3,
        in1(1) => S4602,
        out1 => S5948
    );
nand_n_367: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5948,
        in1(1) => S5943,
        out1 => S5949
    );
nand_n_368: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5949,
        in1(1) => new_datapath_muxmem_in2_3,
        out1 => S5950
    );
notg_369: ENTITY WORK.notg
    PORT MAP (
        in1 => S5950,
        out1 => S5951
    );
nor_n_370: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5949,
        in1(1) => new_datapath_muxmem_in2_3,
        out1 => S5952
    );
nand_n_371: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4289,
        in1(1) => new_controller_fib_2,
        out1 => S5953
    );
nand_n_372: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5903,
        in1(1) => new_controller_outflag_2,
        out1 => S5954
    );
notg_373: ENTITY WORK.notg
    PORT MAP (
        in1 => S5954,
        out1 => S5955
    );
nor_n_374: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5903,
        in1(1) => S3171,
        out1 => S5956
    );
nor_n_375: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5956,
        in1(1) => S5955,
        out1 => S5957
    );
notg_376: ENTITY WORK.notg
    PORT MAP (
        in1 => S5957,
        out1 => new_datapath_addsubunit_in1_2
    );
nand_n_377: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_2,
        in1(1) => S4602,
        out1 => S5958
    );
nand_n_378: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5958,
        in1(1) => S5953,
        out1 => S5959
    );
nand_n_379: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5959,
        in1(1) => new_datapath_muxmem_in2_2,
        out1 => S5960
    );
notg_380: ENTITY WORK.notg
    PORT MAP (
        in1 => S5960,
        out1 => S5961
    );
nand_n_381: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4289,
        in1(1) => new_controller_fib_1,
        out1 => S5962
    );
nand_n_382: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5903,
        in1(1) => new_controller_outflag_1,
        out1 => S5963
    );
notg_383: ENTITY WORK.notg
    PORT MAP (
        in1 => S5963,
        out1 => S5964
    );
nor_n_384: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5903,
        in1(1) => S3160,
        out1 => S5965
    );
nor_n_385: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5965,
        in1(1) => S5964,
        out1 => S5966
    );
notg_386: ENTITY WORK.notg
    PORT MAP (
        in1 => S5966,
        out1 => new_datapath_addsubunit_in1_1
    );
nand_n_387: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_1,
        in1(1) => S4602,
        out1 => S5967
    );
nand_n_388: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5967,
        in1(1) => S5962,
        out1 => S5968
    );
nand_n_389: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5968,
        in1(1) => new_datapath_muxmem_in2_1,
        out1 => S5969
    );
notg_390: ENTITY WORK.notg
    PORT MAP (
        in1 => S5969,
        out1 => S5970
    );
nand_n_391: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4289,
        in1(1) => new_controller_fib_0,
        out1 => S5971
    );
nand_n_392: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5903,
        in1(1) => new_controller_outflag_0,
        out1 => S5972
    );
notg_393: ENTITY WORK.notg
    PORT MAP (
        in1 => S5972,
        out1 => S5973
    );
nor_n_394: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5903,
        in1(1) => S3150,
        out1 => S5974
    );
nor_n_395: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5974,
        in1(1) => S5973,
        out1 => S5975
    );
notg_396: ENTITY WORK.notg
    PORT MAP (
        in1 => S5975,
        out1 => new_datapath_addsubunit_in1_0
    );
nand_n_397: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_0,
        in1(1) => S4602,
        out1 => S5976
    );
nand_n_398: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5976,
        in1(1) => S5971,
        out1 => S5977
    );
notg_399: ENTITY WORK.notg
    PORT MAP (
        in1 => S5977,
        out1 => S5978
    );
nor_n_400: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5978,
        in1(1) => S2625,
        out1 => S5979
    );
nor_n_401: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5968,
        in1(1) => new_datapath_muxmem_in2_1,
        out1 => S5980
    );
nor_n_402: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5980,
        in1(1) => S5970,
        out1 => S5981
    );
nand_n_403: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5981,
        in1(1) => S5979,
        out1 => S5982
    );
nand_n_404: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5982,
        in1(1) => S5969,
        out1 => S5983
    );
nor_n_405: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5959,
        in1(1) => new_datapath_muxmem_in2_2,
        out1 => S5984
    );
nor_n_406: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5984,
        in1(1) => S5961,
        out1 => S5985
    );
nand_n_407: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5985,
        in1(1) => S5983,
        out1 => S5986
    );
nand_n_408: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5986,
        in1(1) => S5960,
        out1 => S5987
    );
nor_n_409: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5987,
        in1(1) => S5951,
        out1 => S5988
    );
nor_n_410: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5988,
        in1(1) => S5952,
        out1 => S5989
    );
nand_n_411: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5989,
        in1(1) => S5942,
        out1 => S5990
    );
nand_n_412: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5990,
        in1(1) => S5939,
        out1 => S5991
    );
nor_n_413: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5991,
        in1(1) => S5930,
        out1 => S5992
    );
nor_n_414: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5992,
        in1(1) => S5931,
        out1 => S5993
    );
nand_n_415: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5993,
        in1(1) => S5922,
        out1 => S5994
    );
nand_n_416: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5994,
        in1(1) => S5919,
        out1 => S5995
    );
nor_n_417: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5995,
        in1(1) => S5911,
        out1 => S5996
    );
nor_n_418: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5996,
        in1(1) => S5912,
        out1 => S5997
    );
nand_n_419: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5997,
        in1(1) => S5018,
        out1 => S5998
    );
nand_n_420: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5998,
        in1(1) => S4986,
        out1 => S5999
    );
nor_n_421: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5999,
        in1(1) => S4943,
        out1 => S6000
    );
nor_n_422: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6000,
        in1(1) => S4954,
        out1 => S6001
    );
nand_n_423: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6001,
        in1(1) => S4900,
        out1 => S6002
    );
nand_n_424: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6002,
        in1(1) => S4868,
        out1 => S6003
    );
nor_n_425: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6003,
        in1(1) => S4836,
        out1 => S6004
    );
nor_n_426: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6004,
        in1(1) => S4825,
        out1 => S6005
    );
nand_n_427: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6005,
        in1(1) => S4783,
        out1 => S6006
    );
nand_n_428: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6006,
        in1(1) => S4750,
        out1 => S6007
    );
nor_n_429: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6007,
        in1(1) => S4708,
        out1 => S6008
    );
nor_n_430: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6008,
        in1(1) => S4718,
        out1 => S6009
    );
nand_n_431: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6009,
        in1(1) => S4665,
        out1 => S6010
    );
nand_n_432: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6010,
        in1(1) => S4632,
        out1 => S6011
    );
nand_n_433: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4602,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S6012
    );
nand_n_434: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6012,
        in1(1) => S4300,
        out1 => S6013
    );
nand_n_435: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6013,
        in1(1) => new_datapath_muxmem_in2_15,
        out1 => S6014
    );
notg_436: ENTITY WORK.notg
    PORT MAP (
        in1 => S6014,
        out1 => S6015
    );
nor_n_437: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6013,
        in1(1) => new_datapath_muxmem_in2_15,
        out1 => S6016
    );
nor_n_438: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6016,
        in1(1) => S6015,
        out1 => S6017
    );
nor_n_439: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6017,
        in1(1) => S6011,
        out1 => S6018
    );
nand_n_440: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5082,
        in1(1) => S4586,
        out1 => S6019
    );
notg_441: ENTITY WORK.notg
    PORT MAP (
        in1 => S6019,
        out1 => S6020
    );
nor_n_442: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6020,
        in1(1) => S4254,
        out1 => S6021
    );
nand_n_443: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6017,
        in1(1) => S6011,
        out1 => S6022
    );
nor_n_444: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6021,
        in1(1) => S6018,
        out1 => S6023
    );
nand_n_445: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6023,
        in1(1) => S6022,
        out1 => S6024
    );
nor_n_446: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4399,
        in1(1) => new_controller_407_B_0,
        out1 => S6025
    );
nor_n_447: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6025,
        in1(1) => S4443,
        out1 => S6026
    );
nor_n_448: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6026,
        in1(1) => S4344,
        out1 => S6027
    );
nor_n_449: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4487,
        in1(1) => new_controller_407_B_0,
        out1 => S6028
    );
nand_n_450: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4421,
        in1(1) => S4344,
        out1 => S6029
    );
nor_n_451: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6029,
        in1(1) => S2996,
        out1 => S6030
    );
nor_n_452: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6030,
        in1(1) => S6028,
        out1 => S6031
    );
nor_n_453: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5061,
        in1(1) => S3117,
        out1 => S6032
    );
nand_n_454: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4355,
        in1(1) => S4322,
        out1 => S6033
    );
nand_n_455: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6033,
        in1(1) => S3969,
        out1 => S6034
    );
nor_n_456: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6034,
        in1(1) => S6032,
        out1 => S6035
    );
nand_n_457: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6035,
        in1(1) => S6031,
        out1 => S6036
    );
nor_n_458: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6036,
        in1(1) => S6027,
        out1 => S6037
    );
nor_n_459: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6037,
        in1(1) => S3958,
        out1 => S6038
    );
nor_n_460: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6038,
        in1(1) => S3936,
        out1 => S6039
    );
nor_n_461: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6039,
        in1(1) => S3771,
        out1 => S6040
    );
nand_n_462: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4155,
        in1(1) => S3719,
        out1 => S6041
    );
nor_n_463: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6041,
        in1(1) => S6040,
        out1 => S6042
    );
nor_n_464: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2636,
        in1(1) => S2625,
        out1 => S6043
    );
nand_n_465: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_muxmem_in2_1,
        in1(1) => new_datapath_muxmem_in2_0,
        out1 => S6044
    );
nor_n_466: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6044,
        in1(1) => S2647,
        out1 => S6045
    );
nand_n_467: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6043,
        in1(1) => new_datapath_muxmem_in2_2,
        out1 => S6046
    );
nor_n_468: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6046,
        in1(1) => S2658,
        out1 => S6047
    );
nand_n_469: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6045,
        in1(1) => new_datapath_muxmem_in2_3,
        out1 => S6048
    );
nand_n_470: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6047,
        in1(1) => new_datapath_muxmem_in2_4,
        out1 => S6049
    );
notg_471: ENTITY WORK.notg
    PORT MAP (
        in1 => S6049,
        out1 => S6050
    );
nand_n_472: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6050,
        in1(1) => new_datapath_muxmem_in2_5,
        out1 => S6051
    );
notg_473: ENTITY WORK.notg
    PORT MAP (
        in1 => S6051,
        out1 => S6052
    );
nand_n_474: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6052,
        in1(1) => new_datapath_muxmem_in2_6,
        out1 => S6053
    );
notg_475: ENTITY WORK.notg
    PORT MAP (
        in1 => S6053,
        out1 => S6054
    );
nand_n_476: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6054,
        in1(1) => new_datapath_muxmem_in2_7,
        out1 => S6055
    );
notg_477: ENTITY WORK.notg
    PORT MAP (
        in1 => S6055,
        out1 => S6056
    );
nor_n_478: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6055,
        in1(1) => S2712,
        out1 => S6057
    );
nand_n_479: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6056,
        in1(1) => new_datapath_muxmem_in2_8,
        out1 => S6058
    );
nor_n_480: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6058,
        in1(1) => S2723,
        out1 => S6059
    );
nand_n_481: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6057,
        in1(1) => new_datapath_muxmem_in2_9,
        out1 => S6060
    );
nor_n_482: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6060,
        in1(1) => S2734,
        out1 => S6061
    );
nand_n_483: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6059,
        in1(1) => new_datapath_muxmem_in2_10,
        out1 => S6062
    );
nand_n_484: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6061,
        in1(1) => new_datapath_muxmem_in2_11,
        out1 => S6063
    );
notg_485: ENTITY WORK.notg
    PORT MAP (
        in1 => S6063,
        out1 => S6064
    );
nand_n_486: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6064,
        in1(1) => new_datapath_muxmem_in2_12,
        out1 => S6065
    );
notg_487: ENTITY WORK.notg
    PORT MAP (
        in1 => S6065,
        out1 => S6066
    );
nor_n_488: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6065,
        in1(1) => S2767,
        out1 => S6067
    );
nand_n_489: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6066,
        in1(1) => new_datapath_muxmem_in2_13,
        out1 => S6068
    );
nand_n_490: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6067,
        in1(1) => new_datapath_muxmem_in2_14,
        out1 => S6069
    );
notg_491: ENTITY WORK.notg
    PORT MAP (
        in1 => S6069,
        out1 => S6070
    );
nand_n_492: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6069,
        in1(1) => new_datapath_muxmem_in2_15,
        out1 => S6071
    );
nor_n_493: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6069,
        in1(1) => new_datapath_muxmem_in2_15,
        out1 => S6072
    );
notg_494: ENTITY WORK.notg
    PORT MAP (
        in1 => S6072,
        out1 => S6073
    );
nand_n_495: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6073,
        in1(1) => S6071,
        out1 => S6074
    );
notg_496: ENTITY WORK.notg
    PORT MAP (
        in1 => S6074,
        out1 => S6075
    );
nor_n_497: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6075,
        in1(1) => S6042,
        out1 => S6076
    );
nand_n_498: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5072,
        in1(1) => new_controller_234_B_0,
        out1 => S6077
    );
notg_499: ENTITY WORK.notg
    PORT MAP (
        in1 => S6077,
        out1 => S6078
    );
nor_n_500: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6078,
        in1(1) => S5408,
        out1 => S6079
    );
nand_n_501: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6077,
        in1(1) => S5419,
        out1 => S6080
    );
nor_n_502: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6079,
        in1(1) => S6076,
        out1 => S6081
    );
nand_n_503: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6081,
        in1(1) => S6024,
        out1 => S6082
    );
nor_n_504: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6080,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S6083
    );
nor_n_505: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6083,
        in1(1) => S4210,
        out1 => S6084
    );
nand_n_506: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6084,
        in1(1) => S6082,
        out1 => S6085
    );
nand_n_507: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6085,
        in1(1) => S4221,
        out1 => S0
    );
nor_n_508: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4133,
        in1(1) => new_controller_pstate_0,
        out1 => S6086
    );
nor_n_509: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => S2581,
        out1 => S1
    );
nand_n_510: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3139,
        in1(1) => S3128,
        out1 => S6087
    );
notg_511: ENTITY WORK.notg
    PORT MAP (
        in1 => S6087,
        out1 => new_controller_1133_S_0
    );
nand_n_512: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_databusin_15,
        out1 => S6088
    );
nand_n_513: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6087,
        in1(1) => new_controller_opcode_7,
        out1 => S6089
    );
nand_n_514: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6089,
        in1(1) => S6088,
        out1 => S2
    );
nor_n_515: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4246,
        in1(1) => new_controller_opcode_3,
        out1 => S6090
    );
nand_n_516: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4238,
        in1(1) => S3062,
        out1 => S6091
    );
nand_n_517: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6091,
        in1(1) => new_datapath_adr_outreg_15,
        out1 => S6092
    );
nand_n_518: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6090,
        in1(1) => S6013,
        out1 => S6093
    );
nand_n_519: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6093,
        in1(1) => S6092,
        out1 => S4
    );
nand_n_520: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4210,
        in1(1) => new_datapath_muxmem_in2_0,
        out1 => S6094
    );
nand_n_521: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5978,
        in1(1) => S2625,
        out1 => S6095
    );
nor_n_522: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6021,
        in1(1) => S5979,
        out1 => S6096
    );
nand_n_523: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6096,
        in1(1) => S6095,
        out1 => S6097
    );
nor_n_524: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6042,
        in1(1) => new_datapath_muxmem_in2_0,
        out1 => S6098
    );
nor_n_525: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6098,
        in1(1) => S6079,
        out1 => S6099
    );
nand_n_526: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6099,
        in1(1) => S6097,
        out1 => S6100
    );
nor_n_527: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6080,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S6101
    );
nor_n_528: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6101,
        in1(1) => S4210,
        out1 => S6102
    );
nand_n_529: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6102,
        in1(1) => S6100,
        out1 => S6103
    );
nand_n_530: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6103,
        in1(1) => S6094,
        out1 => S5
    );
nand_n_531: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4210,
        in1(1) => new_datapath_muxmem_in2_1,
        out1 => S6104
    );
nor_n_532: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5981,
        in1(1) => S5979,
        out1 => S6105
    );
nor_n_533: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6105,
        in1(1) => S6021,
        out1 => S6106
    );
nand_n_534: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6106,
        in1(1) => S5982,
        out1 => S6107
    );
nor_n_535: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_datapath_muxmem_in2_1,
        in1(1) => new_datapath_muxmem_in2_0,
        out1 => S6108
    );
notg_536: ENTITY WORK.notg
    PORT MAP (
        in1 => S6108,
        out1 => S6109
    );
nor_n_537: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6108,
        in1(1) => S6043,
        out1 => S6110
    );
nand_n_538: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6109,
        in1(1) => S6044,
        out1 => S6111
    );
nor_n_539: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6111,
        in1(1) => S6042,
        out1 => S6112
    );
nor_n_540: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6112,
        in1(1) => S6079,
        out1 => S6113
    );
nand_n_541: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6113,
        in1(1) => S6107,
        out1 => S6114
    );
nor_n_542: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6080,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S6115
    );
nor_n_543: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6115,
        in1(1) => S4210,
        out1 => S6116
    );
nand_n_544: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6116,
        in1(1) => S6114,
        out1 => S6117
    );
nand_n_545: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6117,
        in1(1) => S6104,
        out1 => S6
    );
nand_n_546: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4210,
        in1(1) => new_datapath_muxmem_in2_2,
        out1 => S6118
    );
nor_n_547: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5985,
        in1(1) => S5983,
        out1 => S6119
    );
nor_n_548: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6119,
        in1(1) => S6021,
        out1 => S6120
    );
nand_n_549: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6120,
        in1(1) => S5986,
        out1 => S6121
    );
nor_n_550: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6043,
        in1(1) => new_datapath_muxmem_in2_2,
        out1 => S6122
    );
nand_n_551: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6044,
        in1(1) => S2647,
        out1 => S6123
    );
nor_n_552: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6122,
        in1(1) => S6045,
        out1 => S6124
    );
nand_n_553: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6123,
        in1(1) => S6046,
        out1 => S6125
    );
nor_n_554: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6125,
        in1(1) => S6042,
        out1 => S6126
    );
nor_n_555: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6126,
        in1(1) => S6079,
        out1 => S6127
    );
nand_n_556: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6127,
        in1(1) => S6121,
        out1 => S6128
    );
nor_n_557: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6080,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S6129
    );
nor_n_558: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6129,
        in1(1) => S4210,
        out1 => S6130
    );
nand_n_559: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6130,
        in1(1) => S6128,
        out1 => S6131
    );
nand_n_560: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6131,
        in1(1) => S6118,
        out1 => S7
    );
nand_n_561: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4210,
        in1(1) => new_datapath_muxmem_in2_3,
        out1 => S6132
    );
nor_n_562: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5952,
        in1(1) => S5951,
        out1 => S6133
    );
nand_n_563: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6133,
        in1(1) => S5987,
        out1 => S6134
    );
nor_n_564: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6133,
        in1(1) => S5987,
        out1 => S6135
    );
nor_n_565: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6135,
        in1(1) => S6021,
        out1 => S6136
    );
nand_n_566: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6136,
        in1(1) => S6134,
        out1 => S6137
    );
nor_n_567: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6045,
        in1(1) => new_datapath_muxmem_in2_3,
        out1 => S6138
    );
nand_n_568: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6046,
        in1(1) => S2658,
        out1 => S6139
    );
nor_n_569: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6138,
        in1(1) => S6047,
        out1 => S6140
    );
nand_n_570: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6139,
        in1(1) => S6048,
        out1 => S6141
    );
nor_n_571: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6141,
        in1(1) => S6042,
        out1 => S6142
    );
nor_n_572: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6142,
        in1(1) => S6079,
        out1 => S6143
    );
nand_n_573: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6143,
        in1(1) => S6137,
        out1 => S6144
    );
nor_n_574: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6080,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S6145
    );
nor_n_575: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6145,
        in1(1) => S4210,
        out1 => S6146
    );
nand_n_576: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6146,
        in1(1) => S6144,
        out1 => S6147
    );
nand_n_577: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6147,
        in1(1) => S6132,
        out1 => S8
    );
nand_n_578: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4210,
        in1(1) => new_datapath_muxmem_in2_4,
        out1 => S6148
    );
nor_n_579: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5989,
        in1(1) => S5942,
        out1 => S6149
    );
nor_n_580: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6149,
        in1(1) => S6021,
        out1 => S6150
    );
nand_n_581: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6150,
        in1(1) => S5990,
        out1 => S6151
    );
nand_n_582: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6048,
        in1(1) => S2669,
        out1 => S6152
    );
nand_n_583: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6152,
        in1(1) => S6049,
        out1 => S6153
    );
nor_n_584: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6153,
        in1(1) => S6042,
        out1 => S6154
    );
nor_n_585: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6154,
        in1(1) => S6079,
        out1 => S6155
    );
nand_n_586: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6155,
        in1(1) => S6151,
        out1 => S6156
    );
nor_n_587: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6080,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S6157
    );
nor_n_588: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6157,
        in1(1) => S4210,
        out1 => S6158
    );
nand_n_589: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6158,
        in1(1) => S6156,
        out1 => S6159
    );
nand_n_590: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6159,
        in1(1) => S6148,
        out1 => S9
    );
nand_n_591: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4210,
        in1(1) => new_datapath_muxmem_in2_5,
        out1 => S6160
    );
nor_n_592: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5931,
        in1(1) => S5930,
        out1 => S6161
    );
nand_n_593: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6161,
        in1(1) => S5991,
        out1 => S6162
    );
nor_n_594: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6161,
        in1(1) => S5991,
        out1 => S6163
    );
nor_n_595: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6163,
        in1(1) => S6021,
        out1 => S6164
    );
nand_n_596: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6164,
        in1(1) => S6162,
        out1 => S6165
    );
nand_n_597: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6049,
        in1(1) => S2680,
        out1 => S6166
    );
nand_n_598: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6166,
        in1(1) => S6051,
        out1 => S6167
    );
nor_n_599: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6167,
        in1(1) => S6042,
        out1 => S6168
    );
nor_n_600: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6168,
        in1(1) => S6079,
        out1 => S6169
    );
nand_n_601: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6169,
        in1(1) => S6165,
        out1 => S6170
    );
nor_n_602: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6080,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S6171
    );
nor_n_603: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6171,
        in1(1) => S4210,
        out1 => S6172
    );
nand_n_604: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6172,
        in1(1) => S6170,
        out1 => S6173
    );
nand_n_605: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6173,
        in1(1) => S6160,
        out1 => S10
    );
nand_n_606: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4210,
        in1(1) => new_datapath_muxmem_in2_6,
        out1 => S6174
    );
nor_n_607: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5993,
        in1(1) => S5922,
        out1 => S6175
    );
nor_n_608: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6175,
        in1(1) => S6021,
        out1 => S6176
    );
nand_n_609: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6176,
        in1(1) => S5994,
        out1 => S6177
    );
nand_n_610: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6051,
        in1(1) => S2690,
        out1 => S6178
    );
nand_n_611: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6178,
        in1(1) => S6053,
        out1 => S6179
    );
nor_n_612: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6179,
        in1(1) => S6042,
        out1 => S6180
    );
nor_n_613: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6180,
        in1(1) => S6079,
        out1 => S6181
    );
nand_n_614: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6181,
        in1(1) => S6177,
        out1 => S6182
    );
nor_n_615: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6080,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S6183
    );
nor_n_616: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6183,
        in1(1) => S4210,
        out1 => S6184
    );
nand_n_617: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6184,
        in1(1) => S6182,
        out1 => S6185
    );
nand_n_618: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6185,
        in1(1) => S6174,
        out1 => S11
    );
nand_n_619: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4210,
        in1(1) => new_datapath_muxmem_in2_7,
        out1 => S6186
    );
nor_n_620: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5912,
        in1(1) => S5911,
        out1 => S6187
    );
nand_n_621: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6187,
        in1(1) => S5995,
        out1 => S6188
    );
nor_n_622: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6187,
        in1(1) => S5995,
        out1 => S6189
    );
nor_n_623: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6189,
        in1(1) => S6021,
        out1 => S6190
    );
nand_n_624: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6190,
        in1(1) => S6188,
        out1 => S6191
    );
nand_n_625: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6053,
        in1(1) => S2701,
        out1 => S6192
    );
nand_n_626: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6192,
        in1(1) => S6055,
        out1 => S6193
    );
nor_n_627: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6193,
        in1(1) => S6042,
        out1 => S6194
    );
nor_n_628: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6194,
        in1(1) => S6079,
        out1 => S6195
    );
nand_n_629: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6195,
        in1(1) => S6191,
        out1 => S6196
    );
nor_n_630: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6080,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S6197
    );
nor_n_631: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6197,
        in1(1) => S4210,
        out1 => S6198
    );
nand_n_632: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6198,
        in1(1) => S6196,
        out1 => S6199
    );
nand_n_633: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6199,
        in1(1) => S6186,
        out1 => S12
    );
nand_n_634: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4210,
        in1(1) => new_datapath_muxmem_in2_8,
        out1 => S6200
    );
nor_n_635: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5997,
        in1(1) => S5018,
        out1 => S6201
    );
nor_n_636: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6201,
        in1(1) => S6021,
        out1 => S6202
    );
nand_n_637: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6202,
        in1(1) => S5998,
        out1 => S6203
    );
nand_n_638: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6055,
        in1(1) => S2712,
        out1 => S6204
    );
nand_n_639: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6204,
        in1(1) => S6058,
        out1 => S6205
    );
nor_n_640: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6205,
        in1(1) => S6042,
        out1 => S6206
    );
nor_n_641: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6206,
        in1(1) => S6079,
        out1 => S6207
    );
nand_n_642: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6207,
        in1(1) => S6203,
        out1 => S6208
    );
nor_n_643: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6080,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S6209
    );
nor_n_644: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6209,
        in1(1) => S4210,
        out1 => S6210
    );
nand_n_645: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6210,
        in1(1) => S6208,
        out1 => S6211
    );
nand_n_646: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6211,
        in1(1) => S6200,
        out1 => S13
    );
nand_n_647: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4210,
        in1(1) => new_datapath_muxmem_in2_9,
        out1 => S6212
    );
nor_n_648: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4954,
        in1(1) => S4943,
        out1 => S6213
    );
nand_n_649: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6213,
        in1(1) => S5999,
        out1 => S6214
    );
nor_n_650: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6213,
        in1(1) => S5999,
        out1 => S88
    );
nor_n_651: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S88,
        in1(1) => S6021,
        out1 => S89
    );
nand_n_652: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S89,
        in1(1) => S6214,
        out1 => S90
    );
nor_n_653: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6057,
        in1(1) => new_datapath_muxmem_in2_9,
        out1 => S91
    );
nand_n_654: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6058,
        in1(1) => S2723,
        out1 => S92
    );
nor_n_655: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S91,
        in1(1) => S6059,
        out1 => S93
    );
nand_n_656: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S92,
        in1(1) => S6060,
        out1 => S94
    );
nor_n_657: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S94,
        in1(1) => S6042,
        out1 => S95
    );
nor_n_658: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S95,
        in1(1) => S6079,
        out1 => S96
    );
nand_n_659: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S96,
        in1(1) => S90,
        out1 => S97
    );
nor_n_660: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6080,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S98
    );
nor_n_661: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S98,
        in1(1) => S4210,
        out1 => S99
    );
nand_n_662: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S99,
        in1(1) => S97,
        out1 => S100
    );
nand_n_663: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S100,
        in1(1) => S6212,
        out1 => S14
    );
nand_n_664: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4210,
        in1(1) => new_datapath_muxmem_in2_10,
        out1 => S101
    );
nor_n_665: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6001,
        in1(1) => S4900,
        out1 => S102
    );
nor_n_666: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S102,
        in1(1) => S6021,
        out1 => S103
    );
nand_n_667: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S103,
        in1(1) => S6002,
        out1 => S104
    );
nor_n_668: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6059,
        in1(1) => new_datapath_muxmem_in2_10,
        out1 => S105
    );
nand_n_669: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6060,
        in1(1) => S2734,
        out1 => S106
    );
nor_n_670: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S105,
        in1(1) => S6061,
        out1 => S107
    );
nand_n_671: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S106,
        in1(1) => S6062,
        out1 => S108
    );
nor_n_672: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S108,
        in1(1) => S6042,
        out1 => S109
    );
nor_n_673: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S109,
        in1(1) => S6079,
        out1 => S110
    );
nand_n_674: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S110,
        in1(1) => S104,
        out1 => S111
    );
nor_n_675: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6080,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S112
    );
nor_n_676: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S112,
        in1(1) => S4210,
        out1 => S113
    );
nand_n_677: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S113,
        in1(1) => S111,
        out1 => S114
    );
nand_n_678: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S114,
        in1(1) => S101,
        out1 => S15
    );
nand_n_679: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4210,
        in1(1) => new_datapath_muxmem_in2_11,
        out1 => S115
    );
nor_n_680: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4836,
        in1(1) => S4825,
        out1 => S116
    );
nand_n_681: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S116,
        in1(1) => S6003,
        out1 => S117
    );
nor_n_682: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S116,
        in1(1) => S6003,
        out1 => S118
    );
nor_n_683: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S118,
        in1(1) => S6021,
        out1 => S119
    );
nand_n_684: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S119,
        in1(1) => S117,
        out1 => S120
    );
nand_n_685: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6062,
        in1(1) => S2745,
        out1 => S121
    );
nand_n_686: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S121,
        in1(1) => S6063,
        out1 => S122
    );
nor_n_687: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S122,
        in1(1) => S6042,
        out1 => S123
    );
nor_n_688: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S123,
        in1(1) => S6079,
        out1 => S124
    );
nand_n_689: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S124,
        in1(1) => S120,
        out1 => S125
    );
nor_n_690: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6080,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S126
    );
nor_n_691: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S126,
        in1(1) => S4210,
        out1 => S127
    );
nand_n_692: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S127,
        in1(1) => S125,
        out1 => S128
    );
nand_n_693: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S128,
        in1(1) => S115,
        out1 => S16
    );
nand_n_694: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4210,
        in1(1) => new_datapath_muxmem_in2_12,
        out1 => S129
    );
nor_n_695: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6005,
        in1(1) => S4783,
        out1 => S130
    );
nor_n_696: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S130,
        in1(1) => S6021,
        out1 => S131
    );
nand_n_697: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S131,
        in1(1) => S6006,
        out1 => S132
    );
nand_n_698: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6063,
        in1(1) => S2756,
        out1 => S133
    );
nand_n_699: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S133,
        in1(1) => S6065,
        out1 => S134
    );
nor_n_700: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S134,
        in1(1) => S6042,
        out1 => S135
    );
nor_n_701: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S135,
        in1(1) => S6079,
        out1 => S136
    );
nand_n_702: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S136,
        in1(1) => S132,
        out1 => S137
    );
nor_n_703: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6080,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S138
    );
nor_n_704: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S138,
        in1(1) => S4210,
        out1 => S139
    );
nand_n_705: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S139,
        in1(1) => S137,
        out1 => S140
    );
nand_n_706: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S140,
        in1(1) => S129,
        out1 => S17
    );
nand_n_707: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4210,
        in1(1) => new_datapath_muxmem_in2_13,
        out1 => S141
    );
nor_n_708: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4718,
        in1(1) => S4708,
        out1 => S142
    );
nand_n_709: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S142,
        in1(1) => S6007,
        out1 => S143
    );
nor_n_710: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S142,
        in1(1) => S6007,
        out1 => S144
    );
nor_n_711: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S144,
        in1(1) => S6021,
        out1 => S145
    );
nand_n_712: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S145,
        in1(1) => S143,
        out1 => S146
    );
nand_n_713: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6065,
        in1(1) => S2767,
        out1 => S147
    );
nand_n_714: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S147,
        in1(1) => S6068,
        out1 => S148
    );
nor_n_715: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S148,
        in1(1) => S6042,
        out1 => S149
    );
nor_n_716: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S149,
        in1(1) => S6079,
        out1 => S150
    );
nand_n_717: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S150,
        in1(1) => S146,
        out1 => S151
    );
nor_n_718: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6080,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S152
    );
nor_n_719: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S152,
        in1(1) => S4210,
        out1 => S153
    );
nand_n_720: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S153,
        in1(1) => S151,
        out1 => S154
    );
nand_n_721: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S154,
        in1(1) => S141,
        out1 => S18
    );
nand_n_722: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4210,
        in1(1) => new_datapath_muxmem_in2_14,
        out1 => S155
    );
nor_n_723: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6009,
        in1(1) => S4665,
        out1 => S156
    );
nor_n_724: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S156,
        in1(1) => S6021,
        out1 => S157
    );
nand_n_725: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S157,
        in1(1) => S6010,
        out1 => S158
    );
nor_n_726: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6067,
        in1(1) => new_datapath_muxmem_in2_14,
        out1 => S159
    );
nand_n_727: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6068,
        in1(1) => S2778,
        out1 => S160
    );
nor_n_728: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S159,
        in1(1) => S6070,
        out1 => S161
    );
nand_n_729: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S160,
        in1(1) => S6069,
        out1 => S162
    );
nor_n_730: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S162,
        in1(1) => S6042,
        out1 => S163
    );
nor_n_731: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S163,
        in1(1) => S6079,
        out1 => S164
    );
nand_n_732: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S164,
        in1(1) => S158,
        out1 => S165
    );
nor_n_733: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6080,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S166
    );
nor_n_734: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S166,
        in1(1) => S4210,
        out1 => S167
    );
nand_n_735: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S167,
        in1(1) => S165,
        out1 => S168
    );
nand_n_736: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S168,
        in1(1) => S155,
        out1 => S19
    );
nor_n_737: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5719,
        in1(1) => S3062,
        out1 => S169
    );
nor_n_738: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_controller_opcode_2,
        in1(1) => new_controller_234_B_0,
        out1 => S170
    );
nor_n_739: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4578,
        in1(1) => new_controller_opcode_3,
        out1 => S171
    );
notg_740: ENTITY WORK.notg
    PORT MAP (
        in1 => S171,
        out1 => S172
    );
nor_n_741: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_controller_opcode_3,
        in1(1) => new_controller_opcode_2,
        out1 => S173
    );
nand_n_742: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S173,
        in1(1) => S4570,
        out1 => S174
    );
nor_n_743: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S174,
        in1(1) => new_controller_234_B_0,
        out1 => S175
    );
notg_744: ENTITY WORK.notg
    PORT MAP (
        in1 => S175,
        out1 => S176
    );
nand_n_745: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S175,
        in1(1) => new_datapath_instruction_3,
        out1 => S177
    );
notg_746: ENTITY WORK.notg
    PORT MAP (
        in1 => S177,
        out1 => S178
    );
nor_n_747: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S178,
        in1(1) => S169,
        out1 => S179
    );
notg_748: ENTITY WORK.notg
    PORT MAP (
        in1 => S179,
        out1 => new_datapath_muxrs2_outmux_3
    );
nor_n_749: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5719,
        in1(1) => S3029,
        out1 => S180
    );
nand_n_750: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S175,
        in1(1) => new_datapath_instruction_0,
        out1 => S181
    );
notg_751: ENTITY WORK.notg
    PORT MAP (
        in1 => S181,
        out1 => S182
    );
nor_n_752: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S182,
        in1(1) => S180,
        out1 => S183
    );
notg_753: ENTITY WORK.notg
    PORT MAP (
        in1 => S183,
        out1 => new_datapath_muxrs2_outmux_0
    );
nor_n_754: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S183,
        in1(1) => S179,
        out1 => S184
    );
nand_n_755: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_muxrs2_outmux_0,
        in1(1) => new_datapath_muxrs2_outmux_3,
        out1 => S185
    );
nor_n_756: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5719,
        in1(1) => S3040,
        out1 => S186
    );
nand_n_757: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S175,
        in1(1) => new_datapath_instruction_1,
        out1 => S187
    );
notg_758: ENTITY WORK.notg
    PORT MAP (
        in1 => S187,
        out1 => S188
    );
nor_n_759: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S188,
        in1(1) => S186,
        out1 => S189
    );
notg_760: ENTITY WORK.notg
    PORT MAP (
        in1 => S189,
        out1 => new_datapath_muxrs2_outmux_1
    );
nor_n_761: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5719,
        in1(1) => S3051,
        out1 => S190
    );
nand_n_762: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S175,
        in1(1) => new_datapath_instruction_2,
        out1 => S191
    );
notg_763: ENTITY WORK.notg
    PORT MAP (
        in1 => S191,
        out1 => S192
    );
nor_n_764: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S192,
        in1(1) => S190,
        out1 => S193
    );
notg_765: ENTITY WORK.notg
    PORT MAP (
        in1 => S193,
        out1 => new_datapath_muxrs2_outmux_2
    );
nor_n_766: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S193,
        in1(1) => S189,
        out1 => S194
    );
nand_n_767: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_muxrs2_outmux_2,
        in1(1) => new_datapath_muxrs2_outmux_1,
        out1 => S195
    );
nor_n_768: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S195,
        in1(1) => S185,
        out1 => S196
    );
nand_n_769: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S194,
        in1(1) => S184,
        out1 => S197
    );
nand_n_770: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S196,
        in1(1) => new_controller_outflag_6,
        out1 => S198
    );
notg_771: ENTITY WORK.notg
    PORT MAP (
        in1 => S198,
        out1 => S199
    );
nor_n_772: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S196,
        in1(1) => S3303,
        out1 => S200
    );
notg_773: ENTITY WORK.notg
    PORT MAP (
        in1 => S200,
        out1 => S201
    );
nor_n_774: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S200,
        in1(1) => S199,
        out1 => S202
    );
nand_n_775: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S201,
        in1(1) => S198,
        out1 => S203
    );
nand_n_776: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S196,
        in1(1) => new_controller_407_B_2,
        out1 => S204
    );
notg_777: ENTITY WORK.notg
    PORT MAP (
        in1 => S204,
        out1 => S205
    );
nor_n_778: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S196,
        in1(1) => S3292,
        out1 => S206
    );
notg_779: ENTITY WORK.notg
    PORT MAP (
        in1 => S206,
        out1 => S207
    );
nor_n_780: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S206,
        in1(1) => S205,
        out1 => S208
    );
nand_n_781: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S207,
        in1(1) => S204,
        out1 => S209
    );
nor_n_782: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_datapath_multdivunit_1697_B_14,
        in1(1) => new_datapath_multdivunit_1697_B_15,
        out1 => S210
    );
notg_783: ENTITY WORK.notg
    PORT MAP (
        in1 => S210,
        out1 => S211
    );
nor_n_784: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S211,
        in1(1) => new_datapath_multdivunit_1697_B_13,
        out1 => S212
    );
notg_785: ENTITY WORK.notg
    PORT MAP (
        in1 => S212,
        out1 => S213
    );
nor_n_786: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S213,
        in1(1) => new_datapath_multdivunit_1697_B_12,
        out1 => S214
    );
notg_787: ENTITY WORK.notg
    PORT MAP (
        in1 => S214,
        out1 => S215
    );
nor_n_788: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S215,
        in1(1) => new_datapath_multdivunit_1697_B_11,
        out1 => S216
    );
nand_n_789: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S214,
        in1(1) => S3445,
        out1 => S217
    );
nor_n_790: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S217,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S218
    );
notg_791: ENTITY WORK.notg
    PORT MAP (
        in1 => S218,
        out1 => S219
    );
nor_n_792: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S219,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S220
    );
notg_793: ENTITY WORK.notg
    PORT MAP (
        in1 => S220,
        out1 => S221
    );
nor_n_794: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S221,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S222
    );
notg_795: ENTITY WORK.notg
    PORT MAP (
        in1 => S222,
        out1 => S223
    );
nor_n_796: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S197,
        in1(1) => S2614,
        out1 => S224
    );
nand_n_797: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S196,
        in1(1) => new_controller_outflag_7,
        out1 => S225
    );
nor_n_798: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S196,
        in1(1) => S3314,
        out1 => S226
    );
nand_n_799: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S197,
        in1(1) => new_datapath_p2trf_7,
        out1 => S227
    );
nor_n_800: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S226,
        in1(1) => S224,
        out1 => S228
    );
nand_n_801: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S227,
        in1(1) => S225,
        out1 => S229
    );
nor_n_802: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S229,
        in1(1) => S223,
        out1 => S230
    );
nand_n_803: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S228,
        in1(1) => S222,
        out1 => S231
    );
nor_n_804: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S231,
        in1(1) => S203,
        out1 => S232
    );
nand_n_805: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S230,
        in1(1) => S202,
        out1 => S233
    );
nor_n_806: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S233,
        in1(1) => S209,
        out1 => S234
    );
nand_n_807: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S232,
        in1(1) => S208,
        out1 => S235
    );
nand_n_808: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S196,
        in1(1) => new_controller_407_B_0,
        out1 => S236
    );
notg_809: ENTITY WORK.notg
    PORT MAP (
        in1 => S236,
        out1 => S237
    );
nor_n_810: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S196,
        in1(1) => S3281,
        out1 => S238
    );
notg_811: ENTITY WORK.notg
    PORT MAP (
        in1 => S238,
        out1 => S239
    );
nor_n_812: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S238,
        in1(1) => S237,
        out1 => S240
    );
nand_n_813: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S239,
        in1(1) => S236,
        out1 => S241
    );
nor_n_814: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S241,
        in1(1) => S235,
        out1 => S242
    );
nand_n_815: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S240,
        in1(1) => S234,
        out1 => S243
    );
nand_n_816: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S196,
        in1(1) => new_controller_outflag_3,
        out1 => S244
    );
notg_817: ENTITY WORK.notg
    PORT MAP (
        in1 => S244,
        out1 => S245
    );
nor_n_818: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S196,
        in1(1) => S3270,
        out1 => S246
    );
notg_819: ENTITY WORK.notg
    PORT MAP (
        in1 => S246,
        out1 => S247
    );
nor_n_820: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S246,
        in1(1) => S245,
        out1 => S248
    );
nand_n_821: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S247,
        in1(1) => S244,
        out1 => S249
    );
nor_n_822: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S249,
        in1(1) => S243,
        out1 => S250
    );
nand_n_823: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S248,
        in1(1) => S242,
        out1 => S251
    );
nand_n_824: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S196,
        in1(1) => new_controller_outflag_2,
        out1 => S252
    );
notg_825: ENTITY WORK.notg
    PORT MAP (
        in1 => S252,
        out1 => S253
    );
nor_n_826: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S196,
        in1(1) => S3259,
        out1 => S254
    );
notg_827: ENTITY WORK.notg
    PORT MAP (
        in1 => S254,
        out1 => S255
    );
nor_n_828: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S254,
        in1(1) => S253,
        out1 => S256
    );
nand_n_829: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S255,
        in1(1) => S252,
        out1 => S257
    );
nor_n_830: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => S251,
        out1 => S258
    );
nand_n_831: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S256,
        in1(1) => S250,
        out1 => S259
    );
nand_n_832: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S196,
        in1(1) => new_controller_outflag_1,
        out1 => S260
    );
notg_833: ENTITY WORK.notg
    PORT MAP (
        in1 => S260,
        out1 => S261
    );
nor_n_834: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S196,
        in1(1) => S3248,
        out1 => S262
    );
notg_835: ENTITY WORK.notg
    PORT MAP (
        in1 => S262,
        out1 => S263
    );
nor_n_836: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S262,
        in1(1) => S261,
        out1 => S264
    );
nand_n_837: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S263,
        in1(1) => S260,
        out1 => S265
    );
nand_n_838: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S196,
        in1(1) => new_controller_outflag_0,
        out1 => S266
    );
notg_839: ENTITY WORK.notg
    PORT MAP (
        in1 => S266,
        out1 => S267
    );
nor_n_840: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S196,
        in1(1) => S3237,
        out1 => S268
    );
notg_841: ENTITY WORK.notg
    PORT MAP (
        in1 => S268,
        out1 => S269
    );
nor_n_842: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S268,
        in1(1) => S267,
        out1 => S270
    );
nand_n_843: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S269,
        in1(1) => S266,
        out1 => S271
    );
nor_n_844: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S265,
        in1(1) => S259,
        out1 => S272
    );
nand_n_845: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S264,
        in1(1) => S258,
        out1 => S273
    );
nor_n_846: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S273,
        in1(1) => S270,
        out1 => S274
    );
nand_n_847: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S272,
        in1(1) => S271,
        out1 => S275
    );
nor_n_848: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S274,
        in1(1) => S3401,
        out1 => S276
    );
nand_n_849: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S275,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S277
    );
nor_n_850: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S277,
        in1(1) => S265,
        out1 => S278
    );
nand_n_851: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S276,
        in1(1) => S264,
        out1 => S279
    );
nor_n_852: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S264,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S280
    );
nand_n_853: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S265,
        in1(1) => S3401,
        out1 => S281
    );
nor_n_854: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S280,
        in1(1) => S278,
        out1 => S282
    );
nand_n_855: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S281,
        in1(1) => S279,
        out1 => S283
    );
nor_n_856: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S284
    );
nand_n_857: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => S3390,
        out1 => S285
    );
nor_n_858: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S284,
        in1(1) => S283,
        out1 => S286
    );
nand_n_859: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S285,
        in1(1) => S282,
        out1 => S287
    );
nor_n_860: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S286,
        in1(1) => S278,
        out1 => S288
    );
nand_n_861: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S287,
        in1(1) => S279,
        out1 => S289
    );
nor_n_862: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S288,
        in1(1) => S259,
        out1 => S290
    );
nand_n_863: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S289,
        in1(1) => S258,
        out1 => S291
    );
nor_n_864: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S285,
        in1(1) => S282,
        out1 => S292
    );
nor_n_865: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S292,
        in1(1) => S286,
        out1 => S293
    );
nor_n_866: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => S277,
        out1 => S294
    );
nand_n_867: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S291,
        in1(1) => S276,
        out1 => S295
    );
nand_n_868: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S293,
        in1(1) => S290,
        out1 => S296
    );
notg_869: ENTITY WORK.notg
    PORT MAP (
        in1 => S296,
        out1 => S297
    );
nand_n_870: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S296,
        in1(1) => S295,
        out1 => S298
    );
nor_n_871: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S297,
        in1(1) => S294,
        out1 => S299
    );
nor_n_872: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S291,
        in1(1) => S270,
        out1 => S300
    );
nand_n_873: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S290,
        in1(1) => S271,
        out1 => S301
    );
nor_n_874: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S300,
        in1(1) => S3390,
        out1 => S302
    );
nand_n_875: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S301,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S303
    );
nor_n_876: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S303,
        in1(1) => S265,
        out1 => S304
    );
nand_n_877: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S302,
        in1(1) => S264,
        out1 => S305
    );
nor_n_878: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S302,
        in1(1) => S264,
        out1 => S306
    );
nand_n_879: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S303,
        in1(1) => S265,
        out1 => S307
    );
nor_n_880: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S306,
        in1(1) => S304,
        out1 => S308
    );
nand_n_881: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S307,
        in1(1) => S305,
        out1 => S309
    );
nor_n_882: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S310
    );
nand_n_883: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => S3379,
        out1 => S311
    );
nor_n_884: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S310,
        in1(1) => S309,
        out1 => S312
    );
nand_n_885: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S311,
        in1(1) => S308,
        out1 => S313
    );
nor_n_886: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S312,
        in1(1) => S304,
        out1 => S314
    );
nand_n_887: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S313,
        in1(1) => S305,
        out1 => S315
    );
nand_n_888: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => S250,
        out1 => S316
    );
nor_n_889: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S316,
        in1(1) => S314,
        out1 => S317
    );
nand_n_890: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S314,
        in1(1) => S258,
        out1 => S318
    );
nand_n_891: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S318,
        in1(1) => S298,
        out1 => S319
    );
nor_n_892: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S317,
        in1(1) => S299,
        out1 => S320
    );
nor_n_893: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S319,
        in1(1) => S317,
        out1 => S321
    );
nand_n_894: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S320,
        in1(1) => S318,
        out1 => S322
    );
nor_n_895: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S299,
        in1(1) => S257,
        out1 => S323
    );
nand_n_896: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S298,
        in1(1) => S256,
        out1 => S324
    );
nor_n_897: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S323,
        in1(1) => S315,
        out1 => S325
    );
nand_n_898: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S324,
        in1(1) => S314,
        out1 => S326
    );
nor_n_899: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S256,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S327
    );
nand_n_900: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => S3401,
        out1 => S328
    );
nor_n_901: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S327,
        in1(1) => S251,
        out1 => S329
    );
nand_n_902: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S328,
        in1(1) => S250,
        out1 => S330
    );
nor_n_903: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S330,
        in1(1) => S325,
        out1 => S331
    );
nand_n_904: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S329,
        in1(1) => S326,
        out1 => S332
    );
nand_n_905: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S310,
        in1(1) => S309,
        out1 => S333
    );
nand_n_906: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S333,
        in1(1) => S313,
        out1 => S334
    );
nor_n_907: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S331,
        in1(1) => S303,
        out1 => S335
    );
nand_n_908: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S332,
        in1(1) => S302,
        out1 => S336
    );
nor_n_909: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S334,
        in1(1) => S332,
        out1 => S337
    );
notg_910: ENTITY WORK.notg
    PORT MAP (
        in1 => S337,
        out1 => S338
    );
nand_n_911: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S338,
        in1(1) => S336,
        out1 => S339
    );
nor_n_912: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S337,
        in1(1) => S335,
        out1 => S340
    );
nor_n_913: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S340,
        in1(1) => S257,
        out1 => S341
    );
nand_n_914: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S339,
        in1(1) => S256,
        out1 => S342
    );
nor_n_915: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S339,
        in1(1) => S256,
        out1 => S343
    );
nand_n_916: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S340,
        in1(1) => S257,
        out1 => S344
    );
nor_n_917: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S343,
        in1(1) => S341,
        out1 => S345
    );
nand_n_918: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S344,
        in1(1) => S342,
        out1 => S346
    );
nor_n_919: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S331,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S347
    );
nand_n_920: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S332,
        in1(1) => S3379,
        out1 => S348
    );
nor_n_921: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S349
    );
notg_922: ENTITY WORK.notg
    PORT MAP (
        in1 => S349,
        out1 => S350
    );
nor_n_923: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => S3379,
        out1 => S351
    );
nand_n_924: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S352
    );
nand_n_925: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S352,
        in1(1) => S350,
        out1 => S353
    );
nor_n_926: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S351,
        in1(1) => S349,
        out1 => S354
    );
nor_n_927: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S354,
        in1(1) => S332,
        out1 => S355
    );
nand_n_928: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S353,
        in1(1) => S331,
        out1 => S356
    );
nor_n_929: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S355,
        in1(1) => S347,
        out1 => S357
    );
nand_n_930: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S356,
        in1(1) => S348,
        out1 => S358
    );
nor_n_931: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S358,
        in1(1) => S265,
        out1 => S359
    );
nand_n_932: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S357,
        in1(1) => S264,
        out1 => S360
    );
nor_n_933: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S361
    );
nand_n_934: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => S3368,
        out1 => S362
    );
nor_n_935: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S357,
        in1(1) => S264,
        out1 => S363
    );
nand_n_936: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S358,
        in1(1) => S265,
        out1 => S364
    );
nor_n_937: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S363,
        in1(1) => S359,
        out1 => S365
    );
nand_n_938: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S364,
        in1(1) => S360,
        out1 => S366
    );
nor_n_939: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S366,
        in1(1) => S361,
        out1 => S367
    );
nand_n_940: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S365,
        in1(1) => S362,
        out1 => S368
    );
nor_n_941: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S367,
        in1(1) => S359,
        out1 => S369
    );
nand_n_942: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S368,
        in1(1) => S360,
        out1 => S370
    );
nor_n_943: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S369,
        in1(1) => S346,
        out1 => S371
    );
nand_n_944: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S370,
        in1(1) => S345,
        out1 => S372
    );
nor_n_945: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S371,
        in1(1) => S341,
        out1 => S373
    );
nand_n_946: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S372,
        in1(1) => S342,
        out1 => S374
    );
nor_n_947: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S373,
        in1(1) => S249,
        out1 => S375
    );
nand_n_948: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S374,
        in1(1) => S248,
        out1 => S376
    );
nor_n_949: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S374,
        in1(1) => S248,
        out1 => S377
    );
nand_n_950: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S373,
        in1(1) => S249,
        out1 => S378
    );
nor_n_951: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S377,
        in1(1) => S243,
        out1 => S379
    );
nand_n_952: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S378,
        in1(1) => S242,
        out1 => S380
    );
nor_n_953: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S380,
        in1(1) => S375,
        out1 => S381
    );
nor_n_954: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S381,
        in1(1) => S322,
        out1 => S382
    );
notg_955: ENTITY WORK.notg
    PORT MAP (
        in1 => S382,
        out1 => S383
    );
nor_n_956: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S383,
        in1(1) => S241,
        out1 => S384
    );
nand_n_957: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S382,
        in1(1) => S240,
        out1 => S385
    );
nor_n_958: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S321,
        in1(1) => S240,
        out1 => S386
    );
nand_n_959: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S322,
        in1(1) => S241,
        out1 => S387
    );
nor_n_960: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S386,
        in1(1) => S384,
        out1 => S388
    );
nand_n_961: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S387,
        in1(1) => S385,
        out1 => S389
    );
nor_n_962: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S375,
        in1(1) => S321,
        out1 => S390
    );
nand_n_963: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S376,
        in1(1) => S322,
        out1 => S391
    );
nor_n_964: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S390,
        in1(1) => S380,
        out1 => S392
    );
nand_n_965: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S391,
        in1(1) => S379,
        out1 => S393
    );
nor_n_966: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S370,
        in1(1) => S345,
        out1 => S394
    );
nand_n_967: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S369,
        in1(1) => S346,
        out1 => S395
    );
nor_n_968: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S394,
        in1(1) => S371,
        out1 => S396
    );
nand_n_969: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S395,
        in1(1) => S372,
        out1 => S397
    );
nor_n_970: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S396,
        in1(1) => S393,
        out1 => S398
    );
nand_n_971: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S397,
        in1(1) => S392,
        out1 => S399
    );
nor_n_972: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S392,
        in1(1) => S339,
        out1 => S400
    );
nand_n_973: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S393,
        in1(1) => S340,
        out1 => S401
    );
nor_n_974: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S400,
        in1(1) => S398,
        out1 => S402
    );
nand_n_975: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S401,
        in1(1) => S399,
        out1 => S403
    );
nor_n_976: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S403,
        in1(1) => S249,
        out1 => S404
    );
nand_n_977: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S402,
        in1(1) => S248,
        out1 => S405
    );
nor_n_978: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S402,
        in1(1) => S248,
        out1 => S406
    );
nand_n_979: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S403,
        in1(1) => S249,
        out1 => S407
    );
nor_n_980: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S406,
        in1(1) => S404,
        out1 => S408
    );
nand_n_981: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S407,
        in1(1) => S405,
        out1 => S409
    );
nor_n_982: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S365,
        in1(1) => S362,
        out1 => S410
    );
nand_n_983: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S366,
        in1(1) => S361,
        out1 => S411
    );
nor_n_984: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S410,
        in1(1) => S367,
        out1 => S412
    );
nand_n_985: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S411,
        in1(1) => S368,
        out1 => S413
    );
nor_n_986: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S413,
        in1(1) => S393,
        out1 => S414
    );
nand_n_987: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S412,
        in1(1) => S392,
        out1 => S415
    );
nor_n_988: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S392,
        in1(1) => S358,
        out1 => S416
    );
nand_n_989: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S393,
        in1(1) => S357,
        out1 => S417
    );
nor_n_990: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S416,
        in1(1) => S414,
        out1 => S418
    );
nand_n_991: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S417,
        in1(1) => S415,
        out1 => S419
    );
nor_n_992: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S418,
        in1(1) => S257,
        out1 => S420
    );
nand_n_993: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S419,
        in1(1) => S256,
        out1 => S421
    );
nor_n_994: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S419,
        in1(1) => S256,
        out1 => S422
    );
nand_n_995: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S418,
        in1(1) => S257,
        out1 => S423
    );
nor_n_996: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S422,
        in1(1) => S420,
        out1 => S424
    );
nand_n_997: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S423,
        in1(1) => S421,
        out1 => S425
    );
nor_n_998: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => S3368,
        out1 => S426
    );
nand_n_999: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S427
    );
nor_n_1000: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S426,
        in1(1) => S361,
        out1 => S428
    );
nand_n_1001: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S427,
        in1(1) => S362,
        out1 => S429
    );
nor_n_1002: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S428,
        in1(1) => S393,
        out1 => S430
    );
nand_n_1003: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S429,
        in1(1) => S392,
        out1 => S431
    );
nor_n_1004: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S392,
        in1(1) => S3368,
        out1 => S432
    );
nand_n_1005: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S393,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S433
    );
nor_n_1006: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S432,
        in1(1) => S430,
        out1 => S434
    );
nand_n_1007: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S433,
        in1(1) => S431,
        out1 => S435
    );
nor_n_1008: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S434,
        in1(1) => S265,
        out1 => S436
    );
nand_n_1009: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S435,
        in1(1) => S264,
        out1 => S437
    );
nor_n_1010: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S435,
        in1(1) => S264,
        out1 => S438
    );
nand_n_1011: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S434,
        in1(1) => S265,
        out1 => S439
    );
nor_n_1012: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S438,
        in1(1) => S436,
        out1 => S440
    );
nand_n_1013: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S439,
        in1(1) => S437,
        out1 => S441
    );
nor_n_1014: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S442
    );
nand_n_1015: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => S3357,
        out1 => S443
    );
nor_n_1016: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S442,
        in1(1) => S441,
        out1 => S444
    );
nand_n_1017: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S443,
        in1(1) => S440,
        out1 => S445
    );
nor_n_1018: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S444,
        in1(1) => S436,
        out1 => S446
    );
nand_n_1019: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S445,
        in1(1) => S437,
        out1 => S447
    );
nor_n_1020: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S446,
        in1(1) => S425,
        out1 => S448
    );
nand_n_1021: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S447,
        in1(1) => S424,
        out1 => S449
    );
nor_n_1022: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S448,
        in1(1) => S420,
        out1 => S450
    );
nand_n_1023: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S449,
        in1(1) => S421,
        out1 => S451
    );
nor_n_1024: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S450,
        in1(1) => S409,
        out1 => S452
    );
nand_n_1025: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S451,
        in1(1) => S408,
        out1 => S453
    );
nor_n_1026: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S452,
        in1(1) => S404,
        out1 => S454
    );
nand_n_1027: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S453,
        in1(1) => S405,
        out1 => S455
    );
nor_n_1028: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S454,
        in1(1) => S389,
        out1 => S456
    );
nand_n_1029: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S455,
        in1(1) => S388,
        out1 => S457
    );
nor_n_1030: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S456,
        in1(1) => S384,
        out1 => S458
    );
nand_n_1031: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S457,
        in1(1) => S385,
        out1 => S459
    );
nor_n_1032: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S458,
        in1(1) => S235,
        out1 => S460
    );
nand_n_1033: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S459,
        in1(1) => S234,
        out1 => S461
    );
nand_n_1034: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S461,
        in1(1) => S382,
        out1 => S462
    );
nand_n_1035: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S462,
        in1(1) => S296,
        out1 => S463
    );
notg_1036: ENTITY WORK.notg
    PORT MAP (
        in1 => S463,
        out1 => S464
    );
nor_n_1037: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S451,
        in1(1) => S408,
        out1 => S465
    );
nor_n_1038: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S465,
        in1(1) => S452,
        out1 => S466
    );
nor_n_1039: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S466,
        in1(1) => S461,
        out1 => S467
    );
notg_1040: ENTITY WORK.notg
    PORT MAP (
        in1 => S467,
        out1 => S468
    );
nor_n_1041: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S460,
        in1(1) => S402,
        out1 => S469
    );
nand_n_1042: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S461,
        in1(1) => S403,
        out1 => S470
    );
nor_n_1043: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S469,
        in1(1) => S467,
        out1 => S471
    );
nand_n_1044: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S470,
        in1(1) => S468,
        out1 => S472
    );
nor_n_1045: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S472,
        in1(1) => S241,
        out1 => S473
    );
nand_n_1046: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S471,
        in1(1) => S240,
        out1 => S474
    );
nor_n_1047: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S471,
        in1(1) => S240,
        out1 => S475
    );
nand_n_1048: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S472,
        in1(1) => S241,
        out1 => S476
    );
nor_n_1049: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S475,
        in1(1) => S473,
        out1 => S477
    );
nand_n_1050: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S476,
        in1(1) => S474,
        out1 => S478
    );
nor_n_1051: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S447,
        in1(1) => S424,
        out1 => S479
    );
nor_n_1052: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S479,
        in1(1) => S448,
        out1 => S480
    );
nor_n_1053: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S480,
        in1(1) => S461,
        out1 => S481
    );
notg_1054: ENTITY WORK.notg
    PORT MAP (
        in1 => S481,
        out1 => S482
    );
nor_n_1055: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S460,
        in1(1) => S419,
        out1 => S483
    );
nand_n_1056: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S461,
        in1(1) => S418,
        out1 => S484
    );
nor_n_1057: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S483,
        in1(1) => S481,
        out1 => S485
    );
nand_n_1058: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S484,
        in1(1) => S482,
        out1 => S486
    );
nor_n_1059: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S486,
        in1(1) => S249,
        out1 => S487
    );
nand_n_1060: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S485,
        in1(1) => S248,
        out1 => S488
    );
nor_n_1061: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S485,
        in1(1) => S248,
        out1 => S489
    );
nand_n_1062: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S486,
        in1(1) => S249,
        out1 => S490
    );
nor_n_1063: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S489,
        in1(1) => S487,
        out1 => S491
    );
nand_n_1064: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S490,
        in1(1) => S488,
        out1 => S492
    );
nand_n_1065: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S442,
        in1(1) => S441,
        out1 => S493
    );
nand_n_1066: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S493,
        in1(1) => S445,
        out1 => S494
    );
nor_n_1067: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S494,
        in1(1) => S461,
        out1 => S495
    );
notg_1068: ENTITY WORK.notg
    PORT MAP (
        in1 => S495,
        out1 => S496
    );
nand_n_1069: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S461,
        in1(1) => S435,
        out1 => S497
    );
notg_1070: ENTITY WORK.notg
    PORT MAP (
        in1 => S497,
        out1 => S498
    );
nor_n_1071: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S498,
        in1(1) => S495,
        out1 => S499
    );
nand_n_1072: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S497,
        in1(1) => S496,
        out1 => S500
    );
nor_n_1073: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S499,
        in1(1) => S257,
        out1 => S501
    );
nand_n_1074: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S500,
        in1(1) => S256,
        out1 => S502
    );
nor_n_1075: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S500,
        in1(1) => S256,
        out1 => S503
    );
nand_n_1076: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S499,
        in1(1) => S257,
        out1 => S504
    );
nor_n_1077: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S503,
        in1(1) => S501,
        out1 => S505
    );
nand_n_1078: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S504,
        in1(1) => S502,
        out1 => S506
    );
nor_n_1079: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S460,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S507
    );
nand_n_1080: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S461,
        in1(1) => S3357,
        out1 => S508
    );
nor_n_1081: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S509
    );
notg_1082: ENTITY WORK.notg
    PORT MAP (
        in1 => S509,
        out1 => S510
    );
nor_n_1083: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => S3357,
        out1 => S511
    );
nand_n_1084: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S512
    );
nand_n_1085: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S512,
        in1(1) => S510,
        out1 => S513
    );
nor_n_1086: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S511,
        in1(1) => S509,
        out1 => S514
    );
nor_n_1087: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S514,
        in1(1) => S461,
        out1 => S515
    );
nand_n_1088: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S513,
        in1(1) => S460,
        out1 => S516
    );
nor_n_1089: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S515,
        in1(1) => S507,
        out1 => S517
    );
nand_n_1090: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S516,
        in1(1) => S508,
        out1 => S518
    );
nor_n_1091: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S518,
        in1(1) => S265,
        out1 => S519
    );
nand_n_1092: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S517,
        in1(1) => S264,
        out1 => S520
    );
nor_n_1093: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S521
    );
nand_n_1094: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => S3346,
        out1 => S522
    );
nor_n_1095: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S517,
        in1(1) => S264,
        out1 => S523
    );
nand_n_1096: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S518,
        in1(1) => S265,
        out1 => S524
    );
nor_n_1097: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S523,
        in1(1) => S519,
        out1 => S525
    );
nand_n_1098: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S524,
        in1(1) => S520,
        out1 => S526
    );
nor_n_1099: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S526,
        in1(1) => S521,
        out1 => S527
    );
nand_n_1100: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S525,
        in1(1) => S522,
        out1 => S528
    );
nor_n_1101: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S527,
        in1(1) => S519,
        out1 => S529
    );
nand_n_1102: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S528,
        in1(1) => S520,
        out1 => S530
    );
nor_n_1103: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S529,
        in1(1) => S506,
        out1 => S531
    );
nand_n_1104: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S530,
        in1(1) => S505,
        out1 => S532
    );
nor_n_1105: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S531,
        in1(1) => S501,
        out1 => S533
    );
nand_n_1106: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S532,
        in1(1) => S502,
        out1 => S534
    );
nor_n_1107: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S533,
        in1(1) => S492,
        out1 => S535
    );
nand_n_1108: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S534,
        in1(1) => S491,
        out1 => S536
    );
nor_n_1109: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S535,
        in1(1) => S487,
        out1 => S537
    );
nand_n_1110: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S536,
        in1(1) => S488,
        out1 => S538
    );
nor_n_1111: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S537,
        in1(1) => S478,
        out1 => S539
    );
nand_n_1112: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S538,
        in1(1) => S477,
        out1 => S540
    );
nor_n_1113: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S539,
        in1(1) => S473,
        out1 => S541
    );
nand_n_1114: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S540,
        in1(1) => S474,
        out1 => S542
    );
nand_n_1115: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S232,
        in1(1) => S209,
        out1 => S543
    );
nand_n_1116: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S543,
        in1(1) => S542,
        out1 => S544
    );
nand_n_1117: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S541,
        in1(1) => S235,
        out1 => S545
    );
nand_n_1118: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S545,
        in1(1) => S544,
        out1 => S546
    );
nand_n_1119: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S546,
        in1(1) => S463,
        out1 => S547
    );
nor_n_1120: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S464,
        in1(1) => S209,
        out1 => S548
    );
nand_n_1121: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S463,
        in1(1) => S208,
        out1 => S549
    );
nor_n_1122: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S548,
        in1(1) => S542,
        out1 => S550
    );
nand_n_1123: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S549,
        in1(1) => S541,
        out1 => S551
    );
nor_n_1124: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S463,
        in1(1) => S208,
        out1 => S552
    );
nand_n_1125: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S464,
        in1(1) => S209,
        out1 => S553
    );
nor_n_1126: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S552,
        in1(1) => S233,
        out1 => S554
    );
nand_n_1127: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S553,
        in1(1) => S232,
        out1 => S555
    );
nor_n_1128: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S555,
        in1(1) => S550,
        out1 => S556
    );
nand_n_1129: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S554,
        in1(1) => S551,
        out1 => S557
    );
nand_n_1130: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S537,
        in1(1) => S478,
        out1 => S558
    );
nand_n_1131: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S558,
        in1(1) => S540,
        out1 => S559
    );
nand_n_1132: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S559,
        in1(1) => S556,
        out1 => S560
    );
nand_n_1133: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S557,
        in1(1) => S472,
        out1 => S561
    );
nand_n_1134: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S561,
        in1(1) => S560,
        out1 => S562
    );
notg_1135: ENTITY WORK.notg
    PORT MAP (
        in1 => S562,
        out1 => S563
    );
nor_n_1136: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S562,
        in1(1) => S209,
        out1 => S564
    );
nand_n_1137: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S563,
        in1(1) => S208,
        out1 => S565
    );
nor_n_1138: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S563,
        in1(1) => S208,
        out1 => S566
    );
nor_n_1139: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S566,
        in1(1) => S564,
        out1 => S567
    );
notg_1140: ENTITY WORK.notg
    PORT MAP (
        in1 => S567,
        out1 => S568
    );
nand_n_1141: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S533,
        in1(1) => S492,
        out1 => S569
    );
nand_n_1142: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S569,
        in1(1) => S536,
        out1 => S570
    );
nand_n_1143: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S570,
        in1(1) => S556,
        out1 => S571
    );
notg_1144: ENTITY WORK.notg
    PORT MAP (
        in1 => S571,
        out1 => S572
    );
nor_n_1145: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S556,
        in1(1) => S485,
        out1 => S573
    );
notg_1146: ENTITY WORK.notg
    PORT MAP (
        in1 => S573,
        out1 => S574
    );
nor_n_1147: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S573,
        in1(1) => S572,
        out1 => S575
    );
nand_n_1148: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S574,
        in1(1) => S571,
        out1 => S576
    );
nor_n_1149: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S576,
        in1(1) => S241,
        out1 => S577
    );
nand_n_1150: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S575,
        in1(1) => S240,
        out1 => S578
    );
nor_n_1151: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S575,
        in1(1) => S240,
        out1 => S579
    );
nand_n_1152: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S576,
        in1(1) => S241,
        out1 => S580
    );
nor_n_1153: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S579,
        in1(1) => S577,
        out1 => S581
    );
nand_n_1154: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S580,
        in1(1) => S578,
        out1 => S582
    );
nand_n_1155: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S529,
        in1(1) => S506,
        out1 => S583
    );
nand_n_1156: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S583,
        in1(1) => S532,
        out1 => S584
    );
nand_n_1157: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S584,
        in1(1) => S556,
        out1 => S585
    );
nand_n_1158: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S557,
        in1(1) => S499,
        out1 => S586
    );
nand_n_1159: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S586,
        in1(1) => S585,
        out1 => S587
    );
notg_1160: ENTITY WORK.notg
    PORT MAP (
        in1 => S587,
        out1 => S588
    );
nor_n_1161: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S587,
        in1(1) => S249,
        out1 => S589
    );
nand_n_1162: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S588,
        in1(1) => S248,
        out1 => S590
    );
nand_n_1163: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S587,
        in1(1) => S249,
        out1 => S591
    );
notg_1164: ENTITY WORK.notg
    PORT MAP (
        in1 => S591,
        out1 => S592
    );
nor_n_1165: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S592,
        in1(1) => S589,
        out1 => S593
    );
notg_1166: ENTITY WORK.notg
    PORT MAP (
        in1 => S593,
        out1 => S594
    );
nor_n_1167: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S525,
        in1(1) => S522,
        out1 => S595
    );
nand_n_1168: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S526,
        in1(1) => S521,
        out1 => S596
    );
nor_n_1169: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S595,
        in1(1) => S527,
        out1 => S597
    );
nand_n_1170: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S596,
        in1(1) => S528,
        out1 => S598
    );
nor_n_1171: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S598,
        in1(1) => S557,
        out1 => S599
    );
nand_n_1172: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S597,
        in1(1) => S556,
        out1 => S600
    );
nor_n_1173: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S556,
        in1(1) => S518,
        out1 => S601
    );
nand_n_1174: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S557,
        in1(1) => S517,
        out1 => S602
    );
nor_n_1175: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S601,
        in1(1) => S599,
        out1 => S603
    );
nand_n_1176: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S602,
        in1(1) => S600,
        out1 => S604
    );
nor_n_1177: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S603,
        in1(1) => S257,
        out1 => S605
    );
nand_n_1178: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S604,
        in1(1) => S256,
        out1 => S606
    );
nor_n_1179: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S604,
        in1(1) => S256,
        out1 => S607
    );
nand_n_1180: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S603,
        in1(1) => S257,
        out1 => S608
    );
nor_n_1181: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S607,
        in1(1) => S605,
        out1 => S609
    );
nand_n_1182: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S608,
        in1(1) => S606,
        out1 => S610
    );
nor_n_1183: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S556,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S611
    );
nand_n_1184: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S557,
        in1(1) => S3346,
        out1 => S612
    );
nor_n_1185: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => S3346,
        out1 => S613
    );
nand_n_1186: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S614
    );
nor_n_1187: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S613,
        in1(1) => S521,
        out1 => S615
    );
nand_n_1188: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S614,
        in1(1) => S522,
        out1 => S616
    );
nor_n_1189: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S616,
        in1(1) => S557,
        out1 => S617
    );
nand_n_1190: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S615,
        in1(1) => S556,
        out1 => S618
    );
nor_n_1191: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S617,
        in1(1) => S611,
        out1 => S619
    );
nand_n_1192: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S618,
        in1(1) => S612,
        out1 => S620
    );
nor_n_1193: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S620,
        in1(1) => S265,
        out1 => S621
    );
nand_n_1194: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S619,
        in1(1) => S264,
        out1 => S622
    );
nor_n_1195: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S619,
        in1(1) => S264,
        out1 => S623
    );
nand_n_1196: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S620,
        in1(1) => S265,
        out1 => S624
    );
nor_n_1197: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S623,
        in1(1) => S621,
        out1 => S625
    );
nand_n_1198: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S624,
        in1(1) => S622,
        out1 => S626
    );
nor_n_1199: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S627
    );
nand_n_1200: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => S3336,
        out1 => S628
    );
nor_n_1201: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S627,
        in1(1) => S626,
        out1 => S629
    );
nand_n_1202: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S628,
        in1(1) => S625,
        out1 => S630
    );
nor_n_1203: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S629,
        in1(1) => S621,
        out1 => S631
    );
nand_n_1204: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S630,
        in1(1) => S622,
        out1 => S632
    );
nor_n_1205: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S631,
        in1(1) => S610,
        out1 => S633
    );
nand_n_1206: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S632,
        in1(1) => S609,
        out1 => S634
    );
nor_n_1207: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S633,
        in1(1) => S605,
        out1 => S635
    );
nand_n_1208: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S634,
        in1(1) => S606,
        out1 => S636
    );
nor_n_1209: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S635,
        in1(1) => S594,
        out1 => S637
    );
nand_n_1210: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S636,
        in1(1) => S593,
        out1 => S638
    );
nor_n_1211: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S637,
        in1(1) => S589,
        out1 => S639
    );
nand_n_1212: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S638,
        in1(1) => S590,
        out1 => S640
    );
nor_n_1213: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S639,
        in1(1) => S582,
        out1 => S641
    );
nand_n_1214: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S640,
        in1(1) => S581,
        out1 => S642
    );
nor_n_1215: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S641,
        in1(1) => S577,
        out1 => S643
    );
nand_n_1216: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S642,
        in1(1) => S578,
        out1 => S644
    );
nor_n_1217: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S643,
        in1(1) => S568,
        out1 => S645
    );
nand_n_1218: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S644,
        in1(1) => S567,
        out1 => S646
    );
nor_n_1219: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S645,
        in1(1) => S564,
        out1 => S647
    );
nand_n_1220: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S646,
        in1(1) => S565,
        out1 => S648
    );
nand_n_1221: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S230,
        in1(1) => S203,
        out1 => S649
    );
nand_n_1222: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S647,
        in1(1) => S232,
        out1 => S650
    );
nor_n_1223: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S649,
        in1(1) => S647,
        out1 => S651
    );
nor_n_1224: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S651,
        in1(1) => S547,
        out1 => S652
    );
nand_n_1225: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S652,
        in1(1) => S650,
        out1 => S653
    );
notg_1226: ENTITY WORK.notg
    PORT MAP (
        in1 => S653,
        out1 => S654
    );
nor_n_1227: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S547,
        in1(1) => S203,
        out1 => S655
    );
notg_1228: ENTITY WORK.notg
    PORT MAP (
        in1 => S655,
        out1 => S656
    );
nor_n_1229: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S655,
        in1(1) => S648,
        out1 => S657
    );
nand_n_1230: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S656,
        in1(1) => S647,
        out1 => S658
    );
nor_n_1231: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S463,
        in1(1) => S202,
        out1 => S659
    );
nand_n_1232: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S464,
        in1(1) => S203,
        out1 => S660
    );
nor_n_1233: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S659,
        in1(1) => S231,
        out1 => S661
    );
nand_n_1234: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S660,
        in1(1) => S230,
        out1 => S662
    );
nor_n_1235: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S662,
        in1(1) => S657,
        out1 => S663
    );
nand_n_1236: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S661,
        in1(1) => S658,
        out1 => S664
    );
nor_n_1237: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S644,
        in1(1) => S567,
        out1 => S665
    );
nor_n_1238: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S665,
        in1(1) => S645,
        out1 => S666
    );
nor_n_1239: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S666,
        in1(1) => S664,
        out1 => S667
    );
notg_1240: ENTITY WORK.notg
    PORT MAP (
        in1 => S667,
        out1 => S668
    );
nand_n_1241: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S664,
        in1(1) => S562,
        out1 => S669
    );
notg_1242: ENTITY WORK.notg
    PORT MAP (
        in1 => S669,
        out1 => S670
    );
nor_n_1243: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S670,
        in1(1) => S667,
        out1 => S671
    );
nand_n_1244: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S669,
        in1(1) => S668,
        out1 => S672
    );
nor_n_1245: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S672,
        in1(1) => S203,
        out1 => S673
    );
nand_n_1246: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S671,
        in1(1) => S202,
        out1 => S674
    );
nor_n_1247: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S671,
        in1(1) => S202,
        out1 => S675
    );
nand_n_1248: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S672,
        in1(1) => S203,
        out1 => S676
    );
nor_n_1249: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S675,
        in1(1) => S673,
        out1 => S677
    );
nand_n_1250: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S676,
        in1(1) => S674,
        out1 => S678
    );
nand_n_1251: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S639,
        in1(1) => S582,
        out1 => S679
    );
notg_1252: ENTITY WORK.notg
    PORT MAP (
        in1 => S679,
        out1 => S680
    );
nor_n_1253: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S680,
        in1(1) => S641,
        out1 => S681
    );
nor_n_1254: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S681,
        in1(1) => S664,
        out1 => S682
    );
notg_1255: ENTITY WORK.notg
    PORT MAP (
        in1 => S682,
        out1 => S683
    );
nor_n_1256: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S663,
        in1(1) => S575,
        out1 => S684
    );
nand_n_1257: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S664,
        in1(1) => S576,
        out1 => S685
    );
nor_n_1258: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S684,
        in1(1) => S682,
        out1 => S686
    );
nand_n_1259: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S685,
        in1(1) => S683,
        out1 => S687
    );
nor_n_1260: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S687,
        in1(1) => S209,
        out1 => S688
    );
nand_n_1261: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S686,
        in1(1) => S208,
        out1 => S689
    );
nor_n_1262: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S686,
        in1(1) => S208,
        out1 => S690
    );
nand_n_1263: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S687,
        in1(1) => S209,
        out1 => S691
    );
nor_n_1264: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S690,
        in1(1) => S688,
        out1 => S692
    );
nand_n_1265: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S691,
        in1(1) => S689,
        out1 => S693
    );
nand_n_1266: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S635,
        in1(1) => S594,
        out1 => S694
    );
nand_n_1267: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S694,
        in1(1) => S638,
        out1 => S695
    );
nand_n_1268: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S695,
        in1(1) => S663,
        out1 => S696
    );
nand_n_1269: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S664,
        in1(1) => S587,
        out1 => S697
    );
nand_n_1270: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S697,
        in1(1) => S696,
        out1 => S698
    );
notg_1271: ENTITY WORK.notg
    PORT MAP (
        in1 => S698,
        out1 => S699
    );
nor_n_1272: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S698,
        in1(1) => S241,
        out1 => S700
    );
nand_n_1273: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S699,
        in1(1) => S240,
        out1 => S701
    );
nand_n_1274: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S698,
        in1(1) => S241,
        out1 => S702
    );
notg_1275: ENTITY WORK.notg
    PORT MAP (
        in1 => S702,
        out1 => S703
    );
nor_n_1276: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S703,
        in1(1) => S700,
        out1 => S704
    );
notg_1277: ENTITY WORK.notg
    PORT MAP (
        in1 => S704,
        out1 => S705
    );
nand_n_1278: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S631,
        in1(1) => S610,
        out1 => S706
    );
nand_n_1279: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S706,
        in1(1) => S634,
        out1 => S707
    );
nand_n_1280: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S707,
        in1(1) => S663,
        out1 => S708
    );
nand_n_1281: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S664,
        in1(1) => S603,
        out1 => S709
    );
nand_n_1282: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S709,
        in1(1) => S708,
        out1 => S710
    );
notg_1283: ENTITY WORK.notg
    PORT MAP (
        in1 => S710,
        out1 => S711
    );
nor_n_1284: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S710,
        in1(1) => S249,
        out1 => S712
    );
nand_n_1285: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S711,
        in1(1) => S248,
        out1 => S713
    );
nand_n_1286: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S710,
        in1(1) => S249,
        out1 => S714
    );
notg_1287: ENTITY WORK.notg
    PORT MAP (
        in1 => S714,
        out1 => S715
    );
nor_n_1288: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S715,
        in1(1) => S712,
        out1 => S716
    );
notg_1289: ENTITY WORK.notg
    PORT MAP (
        in1 => S716,
        out1 => S717
    );
nor_n_1290: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S628,
        in1(1) => S625,
        out1 => S718
    );
nor_n_1291: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S718,
        in1(1) => S629,
        out1 => S719
    );
nor_n_1292: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S719,
        in1(1) => S664,
        out1 => S720
    );
notg_1293: ENTITY WORK.notg
    PORT MAP (
        in1 => S720,
        out1 => S721
    );
nor_n_1294: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S663,
        in1(1) => S619,
        out1 => S722
    );
nand_n_1295: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S664,
        in1(1) => S620,
        out1 => S723
    );
nor_n_1296: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S722,
        in1(1) => S720,
        out1 => S724
    );
nand_n_1297: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S723,
        in1(1) => S721,
        out1 => S725
    );
nor_n_1298: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S725,
        in1(1) => S257,
        out1 => S726
    );
nand_n_1299: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S724,
        in1(1) => S256,
        out1 => S727
    );
nor_n_1300: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S724,
        in1(1) => S256,
        out1 => S728
    );
nand_n_1301: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S725,
        in1(1) => S257,
        out1 => S729
    );
nor_n_1302: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S728,
        in1(1) => S726,
        out1 => S730
    );
nand_n_1303: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S729,
        in1(1) => S727,
        out1 => S731
    );
nor_n_1304: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S663,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S732
    );
nand_n_1305: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S664,
        in1(1) => S3336,
        out1 => S733
    );
nor_n_1306: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S734
    );
notg_1307: ENTITY WORK.notg
    PORT MAP (
        in1 => S734,
        out1 => S735
    );
nor_n_1308: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => S3336,
        out1 => S736
    );
nand_n_1309: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S737
    );
nand_n_1310: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S737,
        in1(1) => S735,
        out1 => S738
    );
nor_n_1311: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S736,
        in1(1) => S734,
        out1 => S739
    );
nor_n_1312: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S739,
        in1(1) => S664,
        out1 => S740
    );
nand_n_1313: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S738,
        in1(1) => S663,
        out1 => S741
    );
nor_n_1314: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S740,
        in1(1) => S732,
        out1 => S742
    );
nand_n_1315: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S741,
        in1(1) => S733,
        out1 => S743
    );
nor_n_1316: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S743,
        in1(1) => S265,
        out1 => S744
    );
nand_n_1317: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S742,
        in1(1) => S264,
        out1 => S745
    );
nor_n_1318: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S746
    );
nand_n_1319: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => S3325,
        out1 => S747
    );
nor_n_1320: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S742,
        in1(1) => S264,
        out1 => S748
    );
nand_n_1321: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S743,
        in1(1) => S265,
        out1 => S749
    );
nor_n_1322: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S748,
        in1(1) => S744,
        out1 => S750
    );
nand_n_1323: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S749,
        in1(1) => S745,
        out1 => S751
    );
nor_n_1324: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S751,
        in1(1) => S746,
        out1 => S752
    );
nand_n_1325: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S750,
        in1(1) => S747,
        out1 => S753
    );
nor_n_1326: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S752,
        in1(1) => S744,
        out1 => S754
    );
nand_n_1327: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S753,
        in1(1) => S745,
        out1 => S755
    );
nor_n_1328: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S754,
        in1(1) => S731,
        out1 => S756
    );
nand_n_1329: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S755,
        in1(1) => S730,
        out1 => S757
    );
nor_n_1330: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S756,
        in1(1) => S726,
        out1 => S758
    );
nand_n_1331: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S757,
        in1(1) => S727,
        out1 => S759
    );
nor_n_1332: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S758,
        in1(1) => S717,
        out1 => S760
    );
nand_n_1333: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S759,
        in1(1) => S716,
        out1 => S761
    );
nor_n_1334: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S760,
        in1(1) => S712,
        out1 => S762
    );
nand_n_1335: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S761,
        in1(1) => S713,
        out1 => S763
    );
nor_n_1336: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S762,
        in1(1) => S705,
        out1 => S764
    );
nand_n_1337: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S763,
        in1(1) => S704,
        out1 => S765
    );
nor_n_1338: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S764,
        in1(1) => S700,
        out1 => S766
    );
nand_n_1339: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S765,
        in1(1) => S701,
        out1 => S767
    );
nor_n_1340: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S766,
        in1(1) => S693,
        out1 => S768
    );
nand_n_1341: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S767,
        in1(1) => S692,
        out1 => S769
    );
nor_n_1342: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S768,
        in1(1) => S688,
        out1 => S770
    );
nand_n_1343: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S769,
        in1(1) => S689,
        out1 => S771
    );
nor_n_1344: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S770,
        in1(1) => S678,
        out1 => S772
    );
nand_n_1345: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S771,
        in1(1) => S677,
        out1 => S773
    );
nor_n_1346: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S772,
        in1(1) => S673,
        out1 => S774
    );
nand_n_1347: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S773,
        in1(1) => S674,
        out1 => S775
    );
nand_n_1348: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S229,
        in1(1) => S222,
        out1 => S776
    );
nor_n_1349: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S775,
        in1(1) => S231,
        out1 => S777
    );
nor_n_1350: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S776,
        in1(1) => S774,
        out1 => S778
    );
nor_n_1351: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S778,
        in1(1) => S777,
        out1 => S779
    );
nand_n_1352: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S779,
        in1(1) => S654,
        out1 => S780
    );
nand_n_1353: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S547,
        in1(1) => S229,
        out1 => S781
    );
nand_n_1354: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S781,
        in1(1) => S222,
        out1 => S782
    );
notg_1355: ENTITY WORK.notg
    PORT MAP (
        in1 => S782,
        out1 => S783
    );
nor_n_1356: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S782,
        in1(1) => S774,
        out1 => S784
    );
nand_n_1357: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S783,
        in1(1) => S775,
        out1 => S785
    );
nor_n_1358: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S653,
        in1(1) => S231,
        out1 => S786
    );
nand_n_1359: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S654,
        in1(1) => S230,
        out1 => S787
    );
nor_n_1360: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S786,
        in1(1) => S784,
        out1 => S788
    );
nand_n_1361: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S787,
        in1(1) => S785,
        out1 => S789
    );
nand_n_1362: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S770,
        in1(1) => S678,
        out1 => S790
    );
nand_n_1363: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S790,
        in1(1) => S773,
        out1 => S791
    );
nand_n_1364: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S791,
        in1(1) => S789,
        out1 => S792
    );
nand_n_1365: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S788,
        in1(1) => S672,
        out1 => S793
    );
nand_n_1366: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S793,
        in1(1) => S792,
        out1 => S794
    );
notg_1367: ENTITY WORK.notg
    PORT MAP (
        in1 => S794,
        out1 => S795
    );
nor_n_1368: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S794,
        in1(1) => S229,
        out1 => S796
    );
nand_n_1369: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S795,
        in1(1) => S228,
        out1 => S797
    );
nand_n_1370: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S794,
        in1(1) => S229,
        out1 => S798
    );
nand_n_1371: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S798,
        in1(1) => S797,
        out1 => S799
    );
notg_1372: ENTITY WORK.notg
    PORT MAP (
        in1 => S799,
        out1 => S800
    );
nand_n_1373: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S766,
        in1(1) => S693,
        out1 => S801
    );
notg_1374: ENTITY WORK.notg
    PORT MAP (
        in1 => S801,
        out1 => S802
    );
nor_n_1375: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S802,
        in1(1) => S768,
        out1 => S803
    );
nor_n_1376: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S803,
        in1(1) => S788,
        out1 => S804
    );
notg_1377: ENTITY WORK.notg
    PORT MAP (
        in1 => S804,
        out1 => S805
    );
nor_n_1378: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S789,
        in1(1) => S686,
        out1 => S806
    );
nand_n_1379: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S788,
        in1(1) => S687,
        out1 => S807
    );
nor_n_1380: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S806,
        in1(1) => S804,
        out1 => S808
    );
nand_n_1381: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S807,
        in1(1) => S805,
        out1 => S809
    );
nor_n_1382: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S809,
        in1(1) => S203,
        out1 => S810
    );
nand_n_1383: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S808,
        in1(1) => S202,
        out1 => S811
    );
nor_n_1384: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S808,
        in1(1) => S202,
        out1 => S812
    );
nand_n_1385: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S809,
        in1(1) => S203,
        out1 => S813
    );
nor_n_1386: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S763,
        in1(1) => S704,
        out1 => S814
    );
nor_n_1387: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S814,
        in1(1) => S764,
        out1 => S815
    );
nor_n_1388: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S815,
        in1(1) => S788,
        out1 => S816
    );
notg_1389: ENTITY WORK.notg
    PORT MAP (
        in1 => S816,
        out1 => S817
    );
nand_n_1390: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S788,
        in1(1) => S698,
        out1 => S818
    );
notg_1391: ENTITY WORK.notg
    PORT MAP (
        in1 => S818,
        out1 => S819
    );
nor_n_1392: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S819,
        in1(1) => S816,
        out1 => S820
    );
nand_n_1393: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S818,
        in1(1) => S817,
        out1 => S821
    );
nor_n_1394: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S821,
        in1(1) => S209,
        out1 => S822
    );
nand_n_1395: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S820,
        in1(1) => S208,
        out1 => S823
    );
nor_n_1396: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S820,
        in1(1) => S208,
        out1 => S824
    );
nand_n_1397: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S821,
        in1(1) => S209,
        out1 => S825
    );
nor_n_1398: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S824,
        in1(1) => S822,
        out1 => S826
    );
nand_n_1399: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S825,
        in1(1) => S823,
        out1 => S827
    );
nor_n_1400: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S759,
        in1(1) => S716,
        out1 => S828
    );
nor_n_1401: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S828,
        in1(1) => S760,
        out1 => S829
    );
nor_n_1402: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S829,
        in1(1) => S788,
        out1 => S830
    );
notg_1403: ENTITY WORK.notg
    PORT MAP (
        in1 => S830,
        out1 => S831
    );
nand_n_1404: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S788,
        in1(1) => S710,
        out1 => S832
    );
notg_1405: ENTITY WORK.notg
    PORT MAP (
        in1 => S832,
        out1 => S833
    );
nor_n_1406: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S833,
        in1(1) => S830,
        out1 => S834
    );
nand_n_1407: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S832,
        in1(1) => S831,
        out1 => S835
    );
nor_n_1408: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S835,
        in1(1) => S241,
        out1 => S836
    );
nand_n_1409: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S834,
        in1(1) => S240,
        out1 => S837
    );
nor_n_1410: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S834,
        in1(1) => S240,
        out1 => S838
    );
nand_n_1411: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S835,
        in1(1) => S241,
        out1 => S839
    );
nor_n_1412: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S838,
        in1(1) => S836,
        out1 => S840
    );
nand_n_1413: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S839,
        in1(1) => S837,
        out1 => S841
    );
nor_n_1414: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S755,
        in1(1) => S730,
        out1 => S842
    );
nor_n_1415: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S842,
        in1(1) => S756,
        out1 => S843
    );
nor_n_1416: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S843,
        in1(1) => S788,
        out1 => S844
    );
notg_1417: ENTITY WORK.notg
    PORT MAP (
        in1 => S844,
        out1 => S845
    );
nor_n_1418: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S789,
        in1(1) => S724,
        out1 => S846
    );
nand_n_1419: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S788,
        in1(1) => S725,
        out1 => S847
    );
nor_n_1420: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S846,
        in1(1) => S844,
        out1 => S848
    );
nand_n_1421: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S847,
        in1(1) => S845,
        out1 => S849
    );
nor_n_1422: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S849,
        in1(1) => S249,
        out1 => S850
    );
nand_n_1423: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S848,
        in1(1) => S248,
        out1 => S851
    );
nor_n_1424: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S848,
        in1(1) => S248,
        out1 => S852
    );
nand_n_1425: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S849,
        in1(1) => S249,
        out1 => S853
    );
nor_n_1426: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S852,
        in1(1) => S850,
        out1 => S854
    );
nand_n_1427: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S853,
        in1(1) => S851,
        out1 => S855
    );
nor_n_1428: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S750,
        in1(1) => S747,
        out1 => S856
    );
nor_n_1429: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S856,
        in1(1) => S752,
        out1 => S857
    );
nor_n_1430: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S857,
        in1(1) => S788,
        out1 => S858
    );
notg_1431: ENTITY WORK.notg
    PORT MAP (
        in1 => S858,
        out1 => S859
    );
nor_n_1432: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S789,
        in1(1) => S742,
        out1 => S860
    );
nand_n_1433: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S788,
        in1(1) => S743,
        out1 => S861
    );
nor_n_1434: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S860,
        in1(1) => S858,
        out1 => S862
    );
nand_n_1435: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S861,
        in1(1) => S859,
        out1 => S863
    );
nor_n_1436: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S863,
        in1(1) => S257,
        out1 => S864
    );
nand_n_1437: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S862,
        in1(1) => S256,
        out1 => S865
    );
nor_n_1438: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S862,
        in1(1) => S256,
        out1 => S866
    );
nand_n_1439: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S863,
        in1(1) => S257,
        out1 => S867
    );
nor_n_1440: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => S3325,
        out1 => S868
    );
nand_n_1441: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S869
    );
nor_n_1442: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S868,
        in1(1) => S746,
        out1 => S870
    );
nand_n_1443: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S869,
        in1(1) => S747,
        out1 => S871
    );
nor_n_1444: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S871,
        in1(1) => S788,
        out1 => S872
    );
nand_n_1445: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S870,
        in1(1) => S789,
        out1 => S873
    );
nor_n_1446: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S789,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S874
    );
nand_n_1447: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S788,
        in1(1) => S3325,
        out1 => S875
    );
nor_n_1448: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S874,
        in1(1) => S872,
        out1 => S876
    );
nand_n_1449: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S875,
        in1(1) => S873,
        out1 => S877
    );
nor_n_1450: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S877,
        in1(1) => S265,
        out1 => S878
    );
nand_n_1451: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S876,
        in1(1) => S264,
        out1 => S879
    );
nor_n_1452: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S880
    );
nand_n_1453: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => S5916,
        out1 => S881
    );
nor_n_1454: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => S5916,
        out1 => S882
    );
nand_n_1455: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S883
    );
nor_n_1456: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S884
    );
nand_n_1457: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => S5907,
        out1 => S885
    );
nor_n_1458: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => S5907,
        out1 => S886
    );
nand_n_1459: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S887
    );
nor_n_1460: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S886,
        in1(1) => S884,
        out1 => S888
    );
nand_n_1461: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S887,
        in1(1) => S885,
        out1 => S889
    );
nor_n_1462: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S890
    );
nand_n_1463: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => S5907,
        out1 => S891
    );
nor_n_1464: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S876,
        in1(1) => S264,
        out1 => S892
    );
nand_n_1465: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S877,
        in1(1) => S265,
        out1 => S893
    );
nor_n_1466: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S892,
        in1(1) => S878,
        out1 => S894
    );
nand_n_1467: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S893,
        in1(1) => S879,
        out1 => S895
    );
nor_n_1468: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S895,
        in1(1) => S890,
        out1 => S896
    );
nand_n_1469: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S894,
        in1(1) => S891,
        out1 => S897
    );
nor_n_1470: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S896,
        in1(1) => S878,
        out1 => S898
    );
nand_n_1471: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S897,
        in1(1) => S879,
        out1 => S899
    );
nor_n_1472: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S898,
        in1(1) => S866,
        out1 => S900
    );
nand_n_1473: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S899,
        in1(1) => S867,
        out1 => S901
    );
nor_n_1474: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S900,
        in1(1) => S864,
        out1 => S902
    );
nand_n_1475: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S901,
        in1(1) => S865,
        out1 => S903
    );
nor_n_1476: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S902,
        in1(1) => S855,
        out1 => S904
    );
nand_n_1477: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S903,
        in1(1) => S854,
        out1 => S905
    );
nor_n_1478: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S904,
        in1(1) => S850,
        out1 => S906
    );
nand_n_1479: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S905,
        in1(1) => S851,
        out1 => S907
    );
nor_n_1480: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S906,
        in1(1) => S841,
        out1 => S908
    );
nand_n_1481: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S907,
        in1(1) => S840,
        out1 => S909
    );
nor_n_1482: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S908,
        in1(1) => S836,
        out1 => S910
    );
nand_n_1483: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S909,
        in1(1) => S837,
        out1 => S911
    );
nor_n_1484: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S910,
        in1(1) => S827,
        out1 => S912
    );
nand_n_1485: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S911,
        in1(1) => S826,
        out1 => S913
    );
nor_n_1486: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S912,
        in1(1) => S822,
        out1 => S914
    );
nand_n_1487: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S913,
        in1(1) => S823,
        out1 => S915
    );
nor_n_1488: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S914,
        in1(1) => S812,
        out1 => S916
    );
nand_n_1489: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S915,
        in1(1) => S813,
        out1 => S917
    );
nor_n_1490: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S916,
        in1(1) => S810,
        out1 => S918
    );
nand_n_1491: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S917,
        in1(1) => S811,
        out1 => S919
    );
nor_n_1492: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S918,
        in1(1) => S799,
        out1 => S920
    );
nand_n_1493: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S919,
        in1(1) => S800,
        out1 => S921
    );
nor_n_1494: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S920,
        in1(1) => S796,
        out1 => S922
    );
nand_n_1495: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S921,
        in1(1) => S797,
        out1 => S923
    );
nand_n_1496: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S220,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S924
    );
nand_n_1497: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S922,
        in1(1) => S222,
        out1 => S925
    );
nor_n_1498: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S924,
        in1(1) => S922,
        out1 => S926
    );
nor_n_1499: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S926,
        in1(1) => S780,
        out1 => S927
    );
nand_n_1500: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S927,
        in1(1) => S925,
        out1 => S928
    );
nor_n_1501: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S780,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S929
    );
notg_1502: ENTITY WORK.notg
    PORT MAP (
        in1 => S929,
        out1 => S930
    );
nor_n_1503: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S929,
        in1(1) => S923,
        out1 => S931
    );
nand_n_1504: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S930,
        in1(1) => S922,
        out1 => S932
    );
nand_n_1505: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S653,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S933
    );
nand_n_1506: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S933,
        in1(1) => S220,
        out1 => S934
    );
notg_1507: ENTITY WORK.notg
    PORT MAP (
        in1 => S934,
        out1 => S935
    );
nor_n_1508: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S934,
        in1(1) => S931,
        out1 => S936
    );
nand_n_1509: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S935,
        in1(1) => S932,
        out1 => S937
    );
nand_n_1510: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S918,
        in1(1) => S799,
        out1 => S938
    );
nand_n_1511: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S938,
        in1(1) => S921,
        out1 => S939
    );
nand_n_1512: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S939,
        in1(1) => S936,
        out1 => S940
    );
nand_n_1513: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S937,
        in1(1) => S794,
        out1 => S941
    );
nand_n_1514: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S941,
        in1(1) => S940,
        out1 => S942
    );
notg_1515: ENTITY WORK.notg
    PORT MAP (
        in1 => S942,
        out1 => S943
    );
nor_n_1516: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S942,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S944
    );
nand_n_1517: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S943,
        in1(1) => S3478,
        out1 => S945
    );
nand_n_1518: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S942,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S946
    );
notg_1519: ENTITY WORK.notg
    PORT MAP (
        in1 => S946,
        out1 => S947
    );
nor_n_1520: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S947,
        in1(1) => S944,
        out1 => S948
    );
notg_1521: ENTITY WORK.notg
    PORT MAP (
        in1 => S948,
        out1 => S949
    );
nor_n_1522: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S812,
        in1(1) => S810,
        out1 => S950
    );
nand_n_1523: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S813,
        in1(1) => S811,
        out1 => S951
    );
nand_n_1524: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S951,
        in1(1) => S914,
        out1 => S952
    );
nand_n_1525: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S950,
        in1(1) => S915,
        out1 => S953
    );
nand_n_1526: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S953,
        in1(1) => S952,
        out1 => S954
    );
nand_n_1527: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S954,
        in1(1) => S936,
        out1 => S955
    );
nand_n_1528: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S937,
        in1(1) => S809,
        out1 => S956
    );
nand_n_1529: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S956,
        in1(1) => S955,
        out1 => S957
    );
notg_1530: ENTITY WORK.notg
    PORT MAP (
        in1 => S957,
        out1 => S958
    );
nor_n_1531: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S957,
        in1(1) => S229,
        out1 => S959
    );
nand_n_1532: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S958,
        in1(1) => S228,
        out1 => S960
    );
nor_n_1533: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S958,
        in1(1) => S228,
        out1 => S961
    );
nand_n_1534: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S957,
        in1(1) => S229,
        out1 => S962
    );
nor_n_1535: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S911,
        in1(1) => S826,
        out1 => S963
    );
nor_n_1536: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S963,
        in1(1) => S912,
        out1 => S964
    );
nor_n_1537: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S964,
        in1(1) => S937,
        out1 => S965
    );
notg_1538: ENTITY WORK.notg
    PORT MAP (
        in1 => S965,
        out1 => S966
    );
nand_n_1539: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S937,
        in1(1) => S821,
        out1 => S967
    );
notg_1540: ENTITY WORK.notg
    PORT MAP (
        in1 => S967,
        out1 => S968
    );
nor_n_1541: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S968,
        in1(1) => S965,
        out1 => S969
    );
nand_n_1542: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S967,
        in1(1) => S966,
        out1 => S970
    );
nor_n_1543: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S970,
        in1(1) => S203,
        out1 => S971
    );
nand_n_1544: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S969,
        in1(1) => S202,
        out1 => S972
    );
nor_n_1545: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S969,
        in1(1) => S202,
        out1 => S973
    );
nand_n_1546: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S970,
        in1(1) => S203,
        out1 => S974
    );
nor_n_1547: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S973,
        in1(1) => S971,
        out1 => S975
    );
nand_n_1548: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S974,
        in1(1) => S972,
        out1 => S976
    );
nand_n_1549: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S906,
        in1(1) => S841,
        out1 => S977
    );
nand_n_1550: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S977,
        in1(1) => S909,
        out1 => S978
    );
nand_n_1551: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S978,
        in1(1) => S936,
        out1 => S979
    );
nand_n_1552: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S937,
        in1(1) => S835,
        out1 => S980
    );
nand_n_1553: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S980,
        in1(1) => S979,
        out1 => S981
    );
notg_1554: ENTITY WORK.notg
    PORT MAP (
        in1 => S981,
        out1 => S982
    );
nor_n_1555: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S981,
        in1(1) => S209,
        out1 => S983
    );
nand_n_1556: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S982,
        in1(1) => S208,
        out1 => S984
    );
nor_n_1557: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S982,
        in1(1) => S208,
        out1 => S985
    );
nor_n_1558: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S985,
        in1(1) => S983,
        out1 => S986
    );
notg_1559: ENTITY WORK.notg
    PORT MAP (
        in1 => S986,
        out1 => S987
    );
nor_n_1560: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S903,
        in1(1) => S854,
        out1 => S988
    );
nor_n_1561: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S988,
        in1(1) => S904,
        out1 => S989
    );
nor_n_1562: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S989,
        in1(1) => S937,
        out1 => S990
    );
notg_1563: ENTITY WORK.notg
    PORT MAP (
        in1 => S990,
        out1 => S991
    );
nor_n_1564: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S936,
        in1(1) => S848,
        out1 => S992
    );
nand_n_1565: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S937,
        in1(1) => S849,
        out1 => S993
    );
nor_n_1566: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S992,
        in1(1) => S990,
        out1 => S994
    );
nand_n_1567: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S993,
        in1(1) => S991,
        out1 => S995
    );
nor_n_1568: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S995,
        in1(1) => S241,
        out1 => S996
    );
nand_n_1569: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S994,
        in1(1) => S240,
        out1 => S997
    );
nor_n_1570: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S994,
        in1(1) => S240,
        out1 => S998
    );
nand_n_1571: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S995,
        in1(1) => S241,
        out1 => S999
    );
nor_n_1572: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S998,
        in1(1) => S996,
        out1 => S1000
    );
nand_n_1573: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S999,
        in1(1) => S997,
        out1 => S1001
    );
nor_n_1574: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S866,
        in1(1) => S864,
        out1 => S1002
    );
nand_n_1575: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S867,
        in1(1) => S865,
        out1 => S1003
    );
nand_n_1576: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1002,
        in1(1) => S898,
        out1 => S1004
    );
nand_n_1577: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1003,
        in1(1) => S899,
        out1 => S1005
    );
nand_n_1578: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1005,
        in1(1) => S1004,
        out1 => S1006
    );
nor_n_1579: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1006,
        in1(1) => S937,
        out1 => S1007
    );
notg_1580: ENTITY WORK.notg
    PORT MAP (
        in1 => S1007,
        out1 => S1008
    );
nor_n_1581: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S936,
        in1(1) => S862,
        out1 => S1009
    );
nand_n_1582: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S937,
        in1(1) => S863,
        out1 => S1010
    );
nor_n_1583: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1009,
        in1(1) => S1007,
        out1 => S1011
    );
nand_n_1584: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1010,
        in1(1) => S1008,
        out1 => S1012
    );
nor_n_1585: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1012,
        in1(1) => S249,
        out1 => S1013
    );
nor_n_1586: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1011,
        in1(1) => S248,
        out1 => S1014
    );
nor_n_1587: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S894,
        in1(1) => S891,
        out1 => S1015
    );
nor_n_1588: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1015,
        in1(1) => S896,
        out1 => S1016
    );
nor_n_1589: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1016,
        in1(1) => S937,
        out1 => S1017
    );
notg_1590: ENTITY WORK.notg
    PORT MAP (
        in1 => S1017,
        out1 => S1018
    );
nor_n_1591: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S936,
        in1(1) => S876,
        out1 => S1019
    );
nand_n_1592: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S937,
        in1(1) => S877,
        out1 => S1020
    );
nor_n_1593: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1019,
        in1(1) => S1017,
        out1 => S1021
    );
nand_n_1594: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1020,
        in1(1) => S1018,
        out1 => S1022
    );
nor_n_1595: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1022,
        in1(1) => S257,
        out1 => S1023
    );
nand_n_1596: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1021,
        in1(1) => S256,
        out1 => S1024
    );
nor_n_1597: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S937,
        in1(1) => S889,
        out1 => S1025
    );
nand_n_1598: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S936,
        in1(1) => S888,
        out1 => S1026
    );
nor_n_1599: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S936,
        in1(1) => S5907,
        out1 => S1027
    );
nand_n_1600: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S937,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S1028
    );
nor_n_1601: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1027,
        in1(1) => S1025,
        out1 => S1029
    );
nand_n_1602: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1028,
        in1(1) => S1026,
        out1 => S1030
    );
nor_n_1603: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1029,
        in1(1) => S265,
        out1 => S1031
    );
nand_n_1604: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1030,
        in1(1) => S264,
        out1 => S1032
    );
nor_n_1605: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1030,
        in1(1) => S264,
        out1 => S1033
    );
nand_n_1606: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1029,
        in1(1) => S265,
        out1 => S1034
    );
nor_n_1607: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1033,
        in1(1) => S1031,
        out1 => S1035
    );
nand_n_1608: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1034,
        in1(1) => S1032,
        out1 => S1036
    );
nor_n_1609: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1036,
        in1(1) => S880,
        out1 => S1037
    );
nand_n_1610: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1035,
        in1(1) => S881,
        out1 => S1038
    );
nor_n_1611: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1037,
        in1(1) => S1031,
        out1 => S1039
    );
nand_n_1612: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1038,
        in1(1) => S1032,
        out1 => S1040
    );
nor_n_1613: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1021,
        in1(1) => S256,
        out1 => S1041
    );
nor_n_1614: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1041,
        in1(1) => S1023,
        out1 => S1042
    );
notg_1615: ENTITY WORK.notg
    PORT MAP (
        in1 => S1042,
        out1 => S1043
    );
nor_n_1616: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1043,
        in1(1) => S1039,
        out1 => S1044
    );
nand_n_1617: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1042,
        in1(1) => S1040,
        out1 => S1045
    );
nor_n_1618: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1044,
        in1(1) => S1023,
        out1 => S1046
    );
nand_n_1619: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1045,
        in1(1) => S1024,
        out1 => S1047
    );
nor_n_1620: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1046,
        in1(1) => S1014,
        out1 => S1048
    );
nor_n_1621: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1047,
        in1(1) => S1013,
        out1 => S1049
    );
nor_n_1622: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1048,
        in1(1) => S1013,
        out1 => S1050
    );
nor_n_1623: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1049,
        in1(1) => S1014,
        out1 => S1051
    );
nor_n_1624: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1050,
        in1(1) => S1001,
        out1 => S1052
    );
nand_n_1625: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1051,
        in1(1) => S1000,
        out1 => S1053
    );
nor_n_1626: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1052,
        in1(1) => S996,
        out1 => S1054
    );
nand_n_1627: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1053,
        in1(1) => S997,
        out1 => S1055
    );
nor_n_1628: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1054,
        in1(1) => S987,
        out1 => S1056
    );
nand_n_1629: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1055,
        in1(1) => S986,
        out1 => S1057
    );
nor_n_1630: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1056,
        in1(1) => S983,
        out1 => S1058
    );
nand_n_1631: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1057,
        in1(1) => S984,
        out1 => S1059
    );
nor_n_1632: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1058,
        in1(1) => S976,
        out1 => S1060
    );
nand_n_1633: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1059,
        in1(1) => S975,
        out1 => S1061
    );
nor_n_1634: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1060,
        in1(1) => S971,
        out1 => S1062
    );
nand_n_1635: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1061,
        in1(1) => S972,
        out1 => S1063
    );
nor_n_1636: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1062,
        in1(1) => S961,
        out1 => S1064
    );
nand_n_1637: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1063,
        in1(1) => S962,
        out1 => S1065
    );
nor_n_1638: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1064,
        in1(1) => S959,
        out1 => S1066
    );
nand_n_1639: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1065,
        in1(1) => S960,
        out1 => S1067
    );
nor_n_1640: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1066,
        in1(1) => S949,
        out1 => S1068
    );
nand_n_1641: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1067,
        in1(1) => S948,
        out1 => S1069
    );
nor_n_1642: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1068,
        in1(1) => S944,
        out1 => S1070
    );
nand_n_1643: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1069,
        in1(1) => S945,
        out1 => S1071
    );
nand_n_1644: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S218,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S1072
    );
nand_n_1645: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1070,
        in1(1) => S220,
        out1 => S1073
    );
nor_n_1646: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1072,
        in1(1) => S1070,
        out1 => S1074
    );
nor_n_1647: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1074,
        in1(1) => S928,
        out1 => S1075
    );
nand_n_1648: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1075,
        in1(1) => S1073,
        out1 => S1076
    );
nor_n_1649: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S928,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S1077
    );
notg_1650: ENTITY WORK.notg
    PORT MAP (
        in1 => S1077,
        out1 => S1078
    );
nor_n_1651: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1077,
        in1(1) => S1071,
        out1 => S1079
    );
nand_n_1652: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1078,
        in1(1) => S1070,
        out1 => S1080
    );
nand_n_1653: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S780,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S1081
    );
nand_n_1654: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1081,
        in1(1) => S218,
        out1 => S1082
    );
notg_1655: ENTITY WORK.notg
    PORT MAP (
        in1 => S1082,
        out1 => S1083
    );
nor_n_1656: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1082,
        in1(1) => S1079,
        out1 => S1084
    );
nand_n_1657: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1083,
        in1(1) => S1080,
        out1 => S1085
    );
nand_n_1658: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1066,
        in1(1) => S949,
        out1 => S1086
    );
nand_n_1659: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1086,
        in1(1) => S1069,
        out1 => S1087
    );
nand_n_1660: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1087,
        in1(1) => S1084,
        out1 => S1088
    );
nand_n_1661: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1085,
        in1(1) => S942,
        out1 => S1089
    );
nand_n_1662: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1089,
        in1(1) => S1088,
        out1 => S1090
    );
notg_1663: ENTITY WORK.notg
    PORT MAP (
        in1 => S1090,
        out1 => S1091
    );
nor_n_1664: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1090,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S1092
    );
nand_n_1665: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1091,
        in1(1) => S3467,
        out1 => S1093
    );
nand_n_1666: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1090,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S1094
    );
nand_n_1667: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1094,
        in1(1) => S1093,
        out1 => S1095
    );
notg_1668: ENTITY WORK.notg
    PORT MAP (
        in1 => S1095,
        out1 => S1096
    );
nor_n_1669: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S961,
        in1(1) => S959,
        out1 => S1097
    );
nand_n_1670: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S962,
        in1(1) => S960,
        out1 => S1098
    );
nor_n_1671: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1097,
        in1(1) => S1063,
        out1 => S1099
    );
nor_n_1672: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1098,
        in1(1) => S1062,
        out1 => S1100
    );
nor_n_1673: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1100,
        in1(1) => S1099,
        out1 => S1101
    );
nor_n_1674: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1101,
        in1(1) => S1085,
        out1 => S1102
    );
notg_1675: ENTITY WORK.notg
    PORT MAP (
        in1 => S1102,
        out1 => S1103
    );
nand_n_1676: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1085,
        in1(1) => S957,
        out1 => S1104
    );
notg_1677: ENTITY WORK.notg
    PORT MAP (
        in1 => S1104,
        out1 => S1105
    );
nor_n_1678: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1105,
        in1(1) => S1102,
        out1 => S1106
    );
nand_n_1679: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1104,
        in1(1) => S1103,
        out1 => S1107
    );
nor_n_1680: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1107,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S1108
    );
nor_n_1681: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1106,
        in1(1) => S3478,
        out1 => S1109
    );
nand_n_1682: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1058,
        in1(1) => S976,
        out1 => S1110
    );
nand_n_1683: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1110,
        in1(1) => S1061,
        out1 => S1111
    );
nand_n_1684: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1111,
        in1(1) => S1084,
        out1 => S1112
    );
nand_n_1685: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1085,
        in1(1) => S970,
        out1 => S1113
    );
nand_n_1686: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1113,
        in1(1) => S1112,
        out1 => S1114
    );
notg_1687: ENTITY WORK.notg
    PORT MAP (
        in1 => S1114,
        out1 => S1115
    );
nor_n_1688: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1114,
        in1(1) => S229,
        out1 => S1116
    );
nand_n_1689: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1115,
        in1(1) => S228,
        out1 => S1117
    );
nand_n_1690: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1114,
        in1(1) => S229,
        out1 => S1118
    );
nand_n_1691: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1118,
        in1(1) => S1117,
        out1 => S1119
    );
notg_1692: ENTITY WORK.notg
    PORT MAP (
        in1 => S1119,
        out1 => S1120
    );
nor_n_1693: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1055,
        in1(1) => S986,
        out1 => S1121
    );
nor_n_1694: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1121,
        in1(1) => S1056,
        out1 => S1122
    );
nor_n_1695: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1122,
        in1(1) => S1085,
        out1 => S1123
    );
notg_1696: ENTITY WORK.notg
    PORT MAP (
        in1 => S1123,
        out1 => S1124
    );
nand_n_1697: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1085,
        in1(1) => S981,
        out1 => S1125
    );
notg_1698: ENTITY WORK.notg
    PORT MAP (
        in1 => S1125,
        out1 => S1126
    );
nor_n_1699: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1126,
        in1(1) => S1123,
        out1 => S1127
    );
nand_n_1700: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1125,
        in1(1) => S1124,
        out1 => S1128
    );
nor_n_1701: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1128,
        in1(1) => S203,
        out1 => S1129
    );
nand_n_1702: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1127,
        in1(1) => S202,
        out1 => S1130
    );
nor_n_1703: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1127,
        in1(1) => S202,
        out1 => S1131
    );
nand_n_1704: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1128,
        in1(1) => S203,
        out1 => S1132
    );
nor_n_1705: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1131,
        in1(1) => S1129,
        out1 => S1133
    );
nand_n_1706: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1132,
        in1(1) => S1130,
        out1 => S1134
    );
nor_n_1707: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1051,
        in1(1) => S1000,
        out1 => S1135
    );
nor_n_1708: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1135,
        in1(1) => S1052,
        out1 => S1136
    );
nor_n_1709: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1136,
        in1(1) => S1085,
        out1 => S1137
    );
notg_1710: ENTITY WORK.notg
    PORT MAP (
        in1 => S1137,
        out1 => S1138
    );
nor_n_1711: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1084,
        in1(1) => S994,
        out1 => S1139
    );
nand_n_1712: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1085,
        in1(1) => S995,
        out1 => S1140
    );
nor_n_1713: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1139,
        in1(1) => S1137,
        out1 => S1141
    );
nand_n_1714: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1140,
        in1(1) => S1138,
        out1 => S1142
    );
nor_n_1715: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1142,
        in1(1) => S209,
        out1 => S1143
    );
nand_n_1716: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1141,
        in1(1) => S208,
        out1 => S1144
    );
nor_n_1717: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1141,
        in1(1) => S208,
        out1 => S1145
    );
nand_n_1718: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1142,
        in1(1) => S209,
        out1 => S1146
    );
nor_n_1719: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1145,
        in1(1) => S1143,
        out1 => S1147
    );
nand_n_1720: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1146,
        in1(1) => S1144,
        out1 => S1148
    );
nor_n_1721: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1014,
        in1(1) => S1013,
        out1 => S1149
    );
nand_n_1722: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1149,
        in1(1) => S1046,
        out1 => S1150
    );
nor_n_1723: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1149,
        in1(1) => S1046,
        out1 => S1151
    );
notg_1724: ENTITY WORK.notg
    PORT MAP (
        in1 => S1151,
        out1 => S1152
    );
nand_n_1725: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1152,
        in1(1) => S1150,
        out1 => S1153
    );
nor_n_1726: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1153,
        in1(1) => S1085,
        out1 => S1154
    );
notg_1727: ENTITY WORK.notg
    PORT MAP (
        in1 => S1154,
        out1 => S1155
    );
nor_n_1728: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1084,
        in1(1) => S1011,
        out1 => S1156
    );
nand_n_1729: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1085,
        in1(1) => S1012,
        out1 => S1157
    );
nor_n_1730: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1156,
        in1(1) => S1154,
        out1 => S1158
    );
nand_n_1731: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1157,
        in1(1) => S1155,
        out1 => S1159
    );
nor_n_1732: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1159,
        in1(1) => S241,
        out1 => S1160
    );
nand_n_1733: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1158,
        in1(1) => S240,
        out1 => S1161
    );
nor_n_1734: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1158,
        in1(1) => S240,
        out1 => S1162
    );
nand_n_1735: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1159,
        in1(1) => S241,
        out1 => S1163
    );
nor_n_1736: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1162,
        in1(1) => S1160,
        out1 => S1164
    );
nand_n_1737: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1163,
        in1(1) => S1161,
        out1 => S1165
    );
nor_n_1738: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1042,
        in1(1) => S1040,
        out1 => S1166
    );
nor_n_1739: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1166,
        in1(1) => S1044,
        out1 => S1167
    );
nor_n_1740: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1167,
        in1(1) => S1085,
        out1 => S1168
    );
notg_1741: ENTITY WORK.notg
    PORT MAP (
        in1 => S1168,
        out1 => S1169
    );
nand_n_1742: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1085,
        in1(1) => S1022,
        out1 => S1170
    );
notg_1743: ENTITY WORK.notg
    PORT MAP (
        in1 => S1170,
        out1 => S1171
    );
nor_n_1744: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1171,
        in1(1) => S1168,
        out1 => S1172
    );
nand_n_1745: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1170,
        in1(1) => S1169,
        out1 => S1173
    );
nor_n_1746: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1173,
        in1(1) => S249,
        out1 => S1174
    );
nand_n_1747: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1172,
        in1(1) => S248,
        out1 => S1175
    );
nor_n_1748: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1035,
        in1(1) => S881,
        out1 => S1176
    );
nor_n_1749: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1176,
        in1(1) => S1037,
        out1 => S1177
    );
nor_n_1750: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1177,
        in1(1) => S1085,
        out1 => S1178
    );
nor_n_1751: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1084,
        in1(1) => S1030,
        out1 => S1179
    );
nor_n_1752: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1179,
        in1(1) => S1178,
        out1 => S1180
    );
notg_1753: ENTITY WORK.notg
    PORT MAP (
        in1 => S1180,
        out1 => S1181
    );
nor_n_1754: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1181,
        in1(1) => S257,
        out1 => S1182
    );
nand_n_1755: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1180,
        in1(1) => S256,
        out1 => S1183
    );
nor_n_1756: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1180,
        in1(1) => S256,
        out1 => S1184
    );
nand_n_1757: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1181,
        in1(1) => S257,
        out1 => S1185
    );
nor_n_1758: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1184,
        in1(1) => S1182,
        out1 => S1186
    );
nand_n_1759: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1185,
        in1(1) => S1183,
        out1 => S1187
    );
nor_n_1760: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1085,
        in1(1) => S270,
        out1 => S1188
    );
nand_n_1761: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1084,
        in1(1) => S271,
        out1 => S1189
    );
nor_n_1762: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1188,
        in1(1) => S5916,
        out1 => S1190
    );
nand_n_1763: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1189,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S1191
    );
nor_n_1764: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1085,
        in1(1) => S881,
        out1 => S1192
    );
nand_n_1765: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1084,
        in1(1) => S880,
        out1 => S1193
    );
nor_n_1766: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1192,
        in1(1) => S1190,
        out1 => S1194
    );
nand_n_1767: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1193,
        in1(1) => S1191,
        out1 => S1195
    );
nor_n_1768: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1194,
        in1(1) => S265,
        out1 => S1196
    );
nand_n_1769: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1195,
        in1(1) => S264,
        out1 => S1197
    );
nor_n_1770: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1195,
        in1(1) => S264,
        out1 => S1198
    );
nand_n_1771: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1194,
        in1(1) => S265,
        out1 => S1199
    );
nor_n_1772: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1198,
        in1(1) => S1196,
        out1 => S1200
    );
nand_n_1773: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1199,
        in1(1) => S1197,
        out1 => S1201
    );
nor_n_1774: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S1202
    );
nand_n_1775: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => S5936,
        out1 => S1203
    );
nor_n_1776: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => S5936,
        out1 => S1204
    );
nand_n_1777: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S1205
    );
nor_n_1778: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S1206
    );
nand_n_1779: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => S5926,
        out1 => S1207
    );
nor_n_1780: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => S5926,
        out1 => S1208
    );
nand_n_1781: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S1209
    );
nor_n_1782: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1208,
        in1(1) => S1206,
        out1 => S1210
    );
nand_n_1783: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1209,
        in1(1) => S1207,
        out1 => S1211
    );
nor_n_1784: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S1212
    );
nand_n_1785: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => S5926,
        out1 => S1213
    );
nor_n_1786: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1212,
        in1(1) => S1201,
        out1 => S1214
    );
nand_n_1787: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1213,
        in1(1) => S1200,
        out1 => S1215
    );
nor_n_1788: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1214,
        in1(1) => S1196,
        out1 => S1216
    );
nand_n_1789: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1215,
        in1(1) => S1197,
        out1 => S1217
    );
nor_n_1790: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1216,
        in1(1) => S1187,
        out1 => S1218
    );
nand_n_1791: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1217,
        in1(1) => S1186,
        out1 => S1219
    );
nor_n_1792: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1218,
        in1(1) => S1182,
        out1 => S1220
    );
nand_n_1793: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1219,
        in1(1) => S1183,
        out1 => S1221
    );
nor_n_1794: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1172,
        in1(1) => S248,
        out1 => S1222
    );
nand_n_1795: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1173,
        in1(1) => S249,
        out1 => S1223
    );
nor_n_1796: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1222,
        in1(1) => S1174,
        out1 => S1224
    );
nand_n_1797: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1223,
        in1(1) => S1175,
        out1 => S1225
    );
nor_n_1798: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1225,
        in1(1) => S1220,
        out1 => S1226
    );
nand_n_1799: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1224,
        in1(1) => S1221,
        out1 => S1227
    );
nor_n_1800: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1226,
        in1(1) => S1174,
        out1 => S1228
    );
nand_n_1801: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1227,
        in1(1) => S1175,
        out1 => S1229
    );
nor_n_1802: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1228,
        in1(1) => S1165,
        out1 => S1230
    );
nand_n_1803: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1229,
        in1(1) => S1164,
        out1 => S1231
    );
nor_n_1804: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1230,
        in1(1) => S1160,
        out1 => S1232
    );
nand_n_1805: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1231,
        in1(1) => S1161,
        out1 => S1233
    );
nor_n_1806: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1232,
        in1(1) => S1148,
        out1 => S1234
    );
nand_n_1807: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1233,
        in1(1) => S1147,
        out1 => S1235
    );
nor_n_1808: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1234,
        in1(1) => S1143,
        out1 => S1236
    );
nand_n_1809: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1235,
        in1(1) => S1144,
        out1 => S1237
    );
nor_n_1810: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1236,
        in1(1) => S1134,
        out1 => S1238
    );
nand_n_1811: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1237,
        in1(1) => S1133,
        out1 => S1239
    );
nor_n_1812: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1238,
        in1(1) => S1129,
        out1 => S1240
    );
nand_n_1813: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1239,
        in1(1) => S1130,
        out1 => S1241
    );
nor_n_1814: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1240,
        in1(1) => S1119,
        out1 => S1242
    );
nand_n_1815: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1241,
        in1(1) => S1120,
        out1 => S1243
    );
nor_n_1816: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1242,
        in1(1) => S1116,
        out1 => S1244
    );
nand_n_1817: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1243,
        in1(1) => S1117,
        out1 => S1245
    );
nor_n_1818: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1244,
        in1(1) => S1109,
        out1 => S1246
    );
nor_n_1819: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1245,
        in1(1) => S1108,
        out1 => S1247
    );
nor_n_1820: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1246,
        in1(1) => S1108,
        out1 => S1248
    );
nor_n_1821: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1247,
        in1(1) => S1109,
        out1 => S1249
    );
nor_n_1822: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1248,
        in1(1) => S1095,
        out1 => S1250
    );
nand_n_1823: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1249,
        in1(1) => S1096,
        out1 => S1251
    );
nor_n_1824: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1250,
        in1(1) => S1092,
        out1 => S1252
    );
nand_n_1825: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1251,
        in1(1) => S1093,
        out1 => S1253
    );
nand_n_1826: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S216,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S1254
    );
nand_n_1827: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1252,
        in1(1) => S218,
        out1 => S1255
    );
nor_n_1828: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1254,
        in1(1) => S1252,
        out1 => S1256
    );
nor_n_1829: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1256,
        in1(1) => S1076,
        out1 => S1257
    );
nand_n_1830: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1257,
        in1(1) => S1255,
        out1 => S1258
    );
notg_1831: ENTITY WORK.notg
    PORT MAP (
        in1 => S1258,
        out1 => S1259
    );
nor_n_1832: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1076,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S1260
    );
notg_1833: ENTITY WORK.notg
    PORT MAP (
        in1 => S1260,
        out1 => S1261
    );
nor_n_1834: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1260,
        in1(1) => S1253,
        out1 => S1262
    );
nand_n_1835: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1261,
        in1(1) => S1252,
        out1 => S1263
    );
nand_n_1836: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S928,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S1264
    );
nand_n_1837: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1264,
        in1(1) => S216,
        out1 => S1265
    );
notg_1838: ENTITY WORK.notg
    PORT MAP (
        in1 => S1265,
        out1 => S1266
    );
nor_n_1839: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1265,
        in1(1) => S1262,
        out1 => S1267
    );
nand_n_1840: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1266,
        in1(1) => S1263,
        out1 => S1268
    );
nand_n_1841: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1248,
        in1(1) => S1095,
        out1 => S1269
    );
nand_n_1842: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1269,
        in1(1) => S1251,
        out1 => S1270
    );
nand_n_1843: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1270,
        in1(1) => S1267,
        out1 => S1271
    );
nand_n_1844: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1268,
        in1(1) => S1090,
        out1 => S1272
    );
nand_n_1845: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1272,
        in1(1) => S1271,
        out1 => S1273
    );
notg_1846: ENTITY WORK.notg
    PORT MAP (
        in1 => S1273,
        out1 => S1274
    );
nor_n_1847: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1273,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S1275
    );
nand_n_1848: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1274,
        in1(1) => S3456,
        out1 => S1276
    );
nand_n_1849: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1273,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S1277
    );
nand_n_1850: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1277,
        in1(1) => S1276,
        out1 => S1278
    );
notg_1851: ENTITY WORK.notg
    PORT MAP (
        in1 => S1278,
        out1 => S1279
    );
nor_n_1852: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1109,
        in1(1) => S1108,
        out1 => S1280
    );
nor_n_1853: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1280,
        in1(1) => S1245,
        out1 => S1281
    );
nand_n_1854: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1280,
        in1(1) => S1245,
        out1 => S1282
    );
notg_1855: ENTITY WORK.notg
    PORT MAP (
        in1 => S1282,
        out1 => S1283
    );
nor_n_1856: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1283,
        in1(1) => S1281,
        out1 => S1284
    );
nor_n_1857: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1284,
        in1(1) => S1268,
        out1 => S1285
    );
notg_1858: ENTITY WORK.notg
    PORT MAP (
        in1 => S1285,
        out1 => S1286
    );
nand_n_1859: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1268,
        in1(1) => S1107,
        out1 => S1287
    );
notg_1860: ENTITY WORK.notg
    PORT MAP (
        in1 => S1287,
        out1 => S1288
    );
nor_n_1861: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1288,
        in1(1) => S1285,
        out1 => S1289
    );
nand_n_1862: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1287,
        in1(1) => S1286,
        out1 => S1290
    );
nand_n_1863: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1289,
        in1(1) => S3467,
        out1 => S1291
    );
nand_n_1864: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1290,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S1292
    );
nand_n_1865: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1240,
        in1(1) => S1119,
        out1 => S1293
    );
nand_n_1866: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1293,
        in1(1) => S1243,
        out1 => S1294
    );
nand_n_1867: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1294,
        in1(1) => S1267,
        out1 => S1295
    );
nand_n_1868: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1268,
        in1(1) => S1114,
        out1 => S1296
    );
nand_n_1869: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1296,
        in1(1) => S1295,
        out1 => S1297
    );
notg_1870: ENTITY WORK.notg
    PORT MAP (
        in1 => S1297,
        out1 => S1298
    );
nor_n_1871: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1297,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S1299
    );
nand_n_1872: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1298,
        in1(1) => S3478,
        out1 => S1300
    );
nand_n_1873: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1297,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S1301
    );
nand_n_1874: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1301,
        in1(1) => S1300,
        out1 => S1302
    );
notg_1875: ENTITY WORK.notg
    PORT MAP (
        in1 => S1302,
        out1 => S1303
    );
nor_n_1876: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1237,
        in1(1) => S1133,
        out1 => S1304
    );
nor_n_1877: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1304,
        in1(1) => S1238,
        out1 => S1305
    );
nor_n_1878: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1305,
        in1(1) => S1268,
        out1 => S1306
    );
notg_1879: ENTITY WORK.notg
    PORT MAP (
        in1 => S1306,
        out1 => S1307
    );
nand_n_1880: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1268,
        in1(1) => S1128,
        out1 => S1308
    );
notg_1881: ENTITY WORK.notg
    PORT MAP (
        in1 => S1308,
        out1 => S1309
    );
nor_n_1882: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1309,
        in1(1) => S1306,
        out1 => S1310
    );
nand_n_1883: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1308,
        in1(1) => S1307,
        out1 => S1311
    );
nor_n_1884: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1311,
        in1(1) => S229,
        out1 => S1312
    );
nand_n_1885: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1310,
        in1(1) => S228,
        out1 => S1313
    );
nor_n_1886: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1310,
        in1(1) => S228,
        out1 => S1314
    );
nand_n_1887: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1311,
        in1(1) => S229,
        out1 => S1315
    );
nor_n_1888: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1233,
        in1(1) => S1147,
        out1 => S1316
    );
nor_n_1889: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1316,
        in1(1) => S1234,
        out1 => S1317
    );
nor_n_1890: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1317,
        in1(1) => S1268,
        out1 => S1318
    );
notg_1891: ENTITY WORK.notg
    PORT MAP (
        in1 => S1318,
        out1 => S1319
    );
nor_n_1892: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1267,
        in1(1) => S1141,
        out1 => S1320
    );
nand_n_1893: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1268,
        in1(1) => S1142,
        out1 => S1321
    );
nor_n_1894: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1320,
        in1(1) => S1318,
        out1 => S1322
    );
nand_n_1895: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1321,
        in1(1) => S1319,
        out1 => S1323
    );
nor_n_1896: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1323,
        in1(1) => S203,
        out1 => S1324
    );
nand_n_1897: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1322,
        in1(1) => S202,
        out1 => S1325
    );
nor_n_1898: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1322,
        in1(1) => S202,
        out1 => S1326
    );
nand_n_1899: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1323,
        in1(1) => S203,
        out1 => S1327
    );
nor_n_1900: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1326,
        in1(1) => S1324,
        out1 => S1328
    );
nand_n_1901: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1327,
        in1(1) => S1325,
        out1 => S1329
    );
nor_n_1902: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1267,
        in1(1) => S1158,
        out1 => S1330
    );
nand_n_1903: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1268,
        in1(1) => S1159,
        out1 => S1331
    );
nor_n_1904: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1229,
        in1(1) => S1164,
        out1 => S1332
    );
nor_n_1905: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1332,
        in1(1) => S1230,
        out1 => S1333
    );
nor_n_1906: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1333,
        in1(1) => S1268,
        out1 => S1334
    );
notg_1907: ENTITY WORK.notg
    PORT MAP (
        in1 => S1334,
        out1 => S1335
    );
nor_n_1908: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1334,
        in1(1) => S1330,
        out1 => S1336
    );
nand_n_1909: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1335,
        in1(1) => S1331,
        out1 => S1337
    );
nor_n_1910: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1337,
        in1(1) => S209,
        out1 => S1338
    );
nand_n_1911: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1336,
        in1(1) => S208,
        out1 => S1339
    );
nor_n_1912: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1336,
        in1(1) => S208,
        out1 => S1340
    );
nand_n_1913: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1337,
        in1(1) => S209,
        out1 => S1341
    );
nor_n_1914: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1340,
        in1(1) => S1338,
        out1 => S1342
    );
nand_n_1915: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1341,
        in1(1) => S1339,
        out1 => S1343
    );
nand_n_1916: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1268,
        in1(1) => S1173,
        out1 => S1344
    );
notg_1917: ENTITY WORK.notg
    PORT MAP (
        in1 => S1344,
        out1 => S1345
    );
nor_n_1918: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1224,
        in1(1) => S1221,
        out1 => S1346
    );
nor_n_1919: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1346,
        in1(1) => S1226,
        out1 => S1347
    );
nor_n_1920: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1347,
        in1(1) => S1268,
        out1 => S1348
    );
notg_1921: ENTITY WORK.notg
    PORT MAP (
        in1 => S1348,
        out1 => S1349
    );
nor_n_1922: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1348,
        in1(1) => S1345,
        out1 => S1350
    );
nand_n_1923: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1349,
        in1(1) => S1344,
        out1 => S1351
    );
nor_n_1924: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1351,
        in1(1) => S241,
        out1 => S1352
    );
nand_n_1925: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1350,
        in1(1) => S240,
        out1 => S1353
    );
nor_n_1926: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1267,
        in1(1) => S1180,
        out1 => S1354
    );
nand_n_1927: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1268,
        in1(1) => S1181,
        out1 => S1355
    );
nor_n_1928: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1217,
        in1(1) => S1186,
        out1 => S1356
    );
nor_n_1929: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1356,
        in1(1) => S1218,
        out1 => S1357
    );
nor_n_1930: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1357,
        in1(1) => S1268,
        out1 => S1358
    );
notg_1931: ENTITY WORK.notg
    PORT MAP (
        in1 => S1358,
        out1 => S1359
    );
nor_n_1932: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1358,
        in1(1) => S1354,
        out1 => S1360
    );
nand_n_1933: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1359,
        in1(1) => S1355,
        out1 => S1361
    );
nor_n_1934: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1361,
        in1(1) => S249,
        out1 => S1362
    );
nand_n_1935: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1360,
        in1(1) => S248,
        out1 => S1363
    );
nor_n_1936: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1360,
        in1(1) => S248,
        out1 => S1364
    );
nand_n_1937: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1361,
        in1(1) => S249,
        out1 => S1365
    );
nor_n_1938: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1364,
        in1(1) => S1362,
        out1 => S1366
    );
nand_n_1939: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1365,
        in1(1) => S1363,
        out1 => S1367
    );
nor_n_1940: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1213,
        in1(1) => S1200,
        out1 => S1368
    );
nor_n_1941: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1368,
        in1(1) => S1214,
        out1 => S1369
    );
nor_n_1942: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1369,
        in1(1) => S1268,
        out1 => S1370
    );
notg_1943: ENTITY WORK.notg
    PORT MAP (
        in1 => S1370,
        out1 => S1371
    );
nand_n_1944: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1268,
        in1(1) => S1194,
        out1 => S1372
    );
notg_1945: ENTITY WORK.notg
    PORT MAP (
        in1 => S1372,
        out1 => S1373
    );
nor_n_1946: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1373,
        in1(1) => S1370,
        out1 => S1374
    );
nand_n_1947: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1372,
        in1(1) => S1371,
        out1 => S1375
    );
nor_n_1948: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1375,
        in1(1) => S257,
        out1 => S1376
    );
nand_n_1949: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1374,
        in1(1) => S256,
        out1 => S1377
    );
nor_n_1950: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1374,
        in1(1) => S256,
        out1 => S1378
    );
nand_n_1951: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1375,
        in1(1) => S257,
        out1 => S1379
    );
nor_n_1952: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1378,
        in1(1) => S1376,
        out1 => S1380
    );
nand_n_1953: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1379,
        in1(1) => S1377,
        out1 => S1381
    );
nor_n_1954: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1267,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S1382
    );
nand_n_1955: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1268,
        in1(1) => S5926,
        out1 => S1383
    );
nor_n_1956: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1268,
        in1(1) => S1210,
        out1 => S1384
    );
nand_n_1957: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1267,
        in1(1) => S1211,
        out1 => S1385
    );
nor_n_1958: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1384,
        in1(1) => S1382,
        out1 => S1386
    );
nand_n_1959: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1385,
        in1(1) => S1383,
        out1 => S1387
    );
nor_n_1960: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1387,
        in1(1) => S265,
        out1 => S1388
    );
nand_n_1961: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1386,
        in1(1) => S264,
        out1 => S1389
    );
nor_n_1962: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1386,
        in1(1) => S264,
        out1 => S1390
    );
nand_n_1963: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1387,
        in1(1) => S265,
        out1 => S1391
    );
nor_n_1964: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1390,
        in1(1) => S1388,
        out1 => S1392
    );
nand_n_1965: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1391,
        in1(1) => S1389,
        out1 => S1393
    );
nor_n_1966: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1393,
        in1(1) => S1202,
        out1 => S1394
    );
nand_n_1967: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1392,
        in1(1) => S1203,
        out1 => S1395
    );
nor_n_1968: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1394,
        in1(1) => S1388,
        out1 => S1396
    );
nand_n_1969: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1395,
        in1(1) => S1389,
        out1 => S1397
    );
nor_n_1970: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1396,
        in1(1) => S1381,
        out1 => S1398
    );
nand_n_1971: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1397,
        in1(1) => S1380,
        out1 => S1399
    );
nor_n_1972: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1398,
        in1(1) => S1376,
        out1 => S1400
    );
nand_n_1973: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1399,
        in1(1) => S1377,
        out1 => S1401
    );
nor_n_1974: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1400,
        in1(1) => S1367,
        out1 => S1402
    );
nand_n_1975: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1401,
        in1(1) => S1366,
        out1 => S1403
    );
nor_n_1976: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1402,
        in1(1) => S1362,
        out1 => S1404
    );
nand_n_1977: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1403,
        in1(1) => S1363,
        out1 => S1405
    );
nor_n_1978: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1350,
        in1(1) => S240,
        out1 => S1406
    );
nand_n_1979: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1351,
        in1(1) => S241,
        out1 => S1407
    );
nor_n_1980: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1406,
        in1(1) => S1352,
        out1 => S1408
    );
nand_n_1981: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1407,
        in1(1) => S1353,
        out1 => S1409
    );
nor_n_1982: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1409,
        in1(1) => S1404,
        out1 => S1410
    );
nand_n_1983: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1408,
        in1(1) => S1405,
        out1 => S1411
    );
nor_n_1984: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1410,
        in1(1) => S1352,
        out1 => S1412
    );
nand_n_1985: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1411,
        in1(1) => S1353,
        out1 => S1413
    );
nor_n_1986: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1412,
        in1(1) => S1343,
        out1 => S1414
    );
nand_n_1987: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1413,
        in1(1) => S1342,
        out1 => S1415
    );
nor_n_1988: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1414,
        in1(1) => S1338,
        out1 => S1416
    );
nand_n_1989: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1415,
        in1(1) => S1339,
        out1 => S1417
    );
nor_n_1990: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1416,
        in1(1) => S1329,
        out1 => S1418
    );
nand_n_1991: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1417,
        in1(1) => S1328,
        out1 => S1419
    );
nor_n_1992: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1418,
        in1(1) => S1324,
        out1 => S1420
    );
nand_n_1993: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1419,
        in1(1) => S1325,
        out1 => S1421
    );
nor_n_1994: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1420,
        in1(1) => S1314,
        out1 => S1422
    );
nand_n_1995: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1421,
        in1(1) => S1315,
        out1 => S1423
    );
nor_n_1996: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1422,
        in1(1) => S1312,
        out1 => S1424
    );
nand_n_1997: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1423,
        in1(1) => S1313,
        out1 => S1425
    );
nor_n_1998: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1424,
        in1(1) => S1302,
        out1 => S1426
    );
nand_n_1999: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1425,
        in1(1) => S1303,
        out1 => S1427
    );
nor_n_2000: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1426,
        in1(1) => S1299,
        out1 => S1428
    );
nand_n_2001: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1427,
        in1(1) => S1300,
        out1 => S1429
    );
nand_n_2002: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1429,
        in1(1) => S1292,
        out1 => S1430
    );
nand_n_2003: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1428,
        in1(1) => S1291,
        out1 => S1431
    );
nand_n_2004: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1431,
        in1(1) => S1292,
        out1 => S1432
    );
nand_n_2005: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1430,
        in1(1) => S1291,
        out1 => S1433
    );
nor_n_2006: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1432,
        in1(1) => S1278,
        out1 => S1434
    );
nand_n_2007: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1433,
        in1(1) => S1279,
        out1 => S1435
    );
nor_n_2008: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1434,
        in1(1) => S1275,
        out1 => S1436
    );
nand_n_2009: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1435,
        in1(1) => S1276,
        out1 => S1437
    );
nand_n_2010: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S214,
        in1(1) => new_datapath_multdivunit_1697_B_11,
        out1 => S1438
    );
nand_n_2011: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1438,
        in1(1) => S1437,
        out1 => S1439
    );
nand_n_2012: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1436,
        in1(1) => S217,
        out1 => S1440
    );
nand_n_2013: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1440,
        in1(1) => S1439,
        out1 => S1441
    );
nand_n_2014: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1441,
        in1(1) => S1259,
        out1 => S1442
    );
nor_n_2015: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1442,
        in1(1) => new_datapath_multdivunit_1697_B_12,
        out1 => S1443
    );
notg_2016: ENTITY WORK.notg
    PORT MAP (
        in1 => S1443,
        out1 => S1444
    );
nand_n_2017: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1076,
        in1(1) => new_datapath_multdivunit_1697_B_11,
        out1 => S1445
    );
nand_n_2018: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1445,
        in1(1) => S214,
        out1 => S1446
    );
notg_2019: ENTITY WORK.notg
    PORT MAP (
        in1 => S1446,
        out1 => S1447
    );
nor_n_2020: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1446,
        in1(1) => S1436,
        out1 => S1448
    );
nand_n_2021: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1447,
        in1(1) => S1437,
        out1 => S1449
    );
nor_n_2022: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1258,
        in1(1) => S217,
        out1 => S1450
    );
nand_n_2023: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1259,
        in1(1) => S216,
        out1 => S1451
    );
nor_n_2024: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1450,
        in1(1) => S1448,
        out1 => S1452
    );
nand_n_2025: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1451,
        in1(1) => S1449,
        out1 => S1453
    );
nand_n_2026: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1432,
        in1(1) => S1278,
        out1 => S1454
    );
nand_n_2027: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1454,
        in1(1) => S1435,
        out1 => S1455
    );
nand_n_2028: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1455,
        in1(1) => S1453,
        out1 => S1456
    );
nand_n_2029: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1452,
        in1(1) => S1273,
        out1 => S1457
    );
nand_n_2030: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1457,
        in1(1) => S1456,
        out1 => S1458
    );
notg_2031: ENTITY WORK.notg
    PORT MAP (
        in1 => S1458,
        out1 => S1459
    );
nor_n_2032: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1458,
        in1(1) => new_datapath_multdivunit_1697_B_11,
        out1 => S1460
    );
nand_n_2033: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1459,
        in1(1) => S3445,
        out1 => S1461
    );
nand_n_2034: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1458,
        in1(1) => new_datapath_multdivunit_1697_B_11,
        out1 => S1462
    );
nand_n_2035: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1462,
        in1(1) => S1461,
        out1 => S1463
    );
notg_2036: ENTITY WORK.notg
    PORT MAP (
        in1 => S1463,
        out1 => S1464
    );
nand_n_2037: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1292,
        in1(1) => S1291,
        out1 => S1465
    );
nand_n_2038: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1465,
        in1(1) => S1429,
        out1 => S1466
    );
notg_2039: ENTITY WORK.notg
    PORT MAP (
        in1 => S1466,
        out1 => S1467
    );
nor_n_2040: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1465,
        in1(1) => S1429,
        out1 => S1468
    );
nor_n_2041: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1468,
        in1(1) => S1467,
        out1 => S1469
    );
nor_n_2042: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1469,
        in1(1) => S1452,
        out1 => S1470
    );
notg_2043: ENTITY WORK.notg
    PORT MAP (
        in1 => S1470,
        out1 => S1471
    );
nand_n_2044: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1452,
        in1(1) => S1289,
        out1 => S1472
    );
notg_2045: ENTITY WORK.notg
    PORT MAP (
        in1 => S1472,
        out1 => S1473
    );
nor_n_2046: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1473,
        in1(1) => S1470,
        out1 => S1474
    );
nand_n_2047: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1472,
        in1(1) => S1471,
        out1 => S1475
    );
nor_n_2048: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1475,
        in1(1) => S3456,
        out1 => S1476
    );
nor_n_2049: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1474,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S1477
    );
nand_n_2050: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1424,
        in1(1) => S1302,
        out1 => S1478
    );
nand_n_2051: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1478,
        in1(1) => S1427,
        out1 => S1479
    );
nand_n_2052: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1479,
        in1(1) => S1453,
        out1 => S1480
    );
nand_n_2053: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1452,
        in1(1) => S1297,
        out1 => S1481
    );
nand_n_2054: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1481,
        in1(1) => S1480,
        out1 => S1482
    );
notg_2055: ENTITY WORK.notg
    PORT MAP (
        in1 => S1482,
        out1 => S1483
    );
nor_n_2056: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1482,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S1484
    );
nand_n_2057: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1483,
        in1(1) => S3467,
        out1 => S1485
    );
nand_n_2058: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1482,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S1486
    );
nand_n_2059: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1486,
        in1(1) => S1485,
        out1 => S1487
    );
notg_2060: ENTITY WORK.notg
    PORT MAP (
        in1 => S1487,
        out1 => S1488
    );
nor_n_2061: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1314,
        in1(1) => S1312,
        out1 => S1489
    );
nand_n_2062: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1315,
        in1(1) => S1313,
        out1 => S1490
    );
nor_n_2063: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1489,
        in1(1) => S1421,
        out1 => S1491
    );
nor_n_2064: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1490,
        in1(1) => S1420,
        out1 => S1492
    );
nor_n_2065: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1492,
        in1(1) => S1491,
        out1 => S1493
    );
nor_n_2066: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1493,
        in1(1) => S1452,
        out1 => S1494
    );
notg_2067: ENTITY WORK.notg
    PORT MAP (
        in1 => S1494,
        out1 => S1495
    );
nand_n_2068: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1452,
        in1(1) => S1311,
        out1 => S1496
    );
notg_2069: ENTITY WORK.notg
    PORT MAP (
        in1 => S1496,
        out1 => S1497
    );
nor_n_2070: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1497,
        in1(1) => S1494,
        out1 => S1498
    );
nand_n_2071: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1496,
        in1(1) => S1495,
        out1 => S1499
    );
nor_n_2072: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1499,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S1500
    );
nor_n_2073: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1498,
        in1(1) => S3478,
        out1 => S1501
    );
nand_n_2074: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1416,
        in1(1) => S1329,
        out1 => S1502
    );
nand_n_2075: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1502,
        in1(1) => S1419,
        out1 => S1503
    );
nand_n_2076: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1503,
        in1(1) => S1453,
        out1 => S1504
    );
nand_n_2077: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1452,
        in1(1) => S1323,
        out1 => S1505
    );
nand_n_2078: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1505,
        in1(1) => S1504,
        out1 => S1506
    );
notg_2079: ENTITY WORK.notg
    PORT MAP (
        in1 => S1506,
        out1 => S1507
    );
nor_n_2080: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1506,
        in1(1) => S229,
        out1 => S1508
    );
nand_n_2081: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1507,
        in1(1) => S228,
        out1 => S1509
    );
nand_n_2082: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1506,
        in1(1) => S229,
        out1 => S1510
    );
nand_n_2083: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1510,
        in1(1) => S1509,
        out1 => S1511
    );
notg_2084: ENTITY WORK.notg
    PORT MAP (
        in1 => S1511,
        out1 => S1512
    );
nor_n_2085: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1413,
        in1(1) => S1342,
        out1 => S1513
    );
nor_n_2086: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1513,
        in1(1) => S1414,
        out1 => S1514
    );
nor_n_2087: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1514,
        in1(1) => S1452,
        out1 => S1515
    );
notg_2088: ENTITY WORK.notg
    PORT MAP (
        in1 => S1515,
        out1 => S1516
    );
nand_n_2089: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1452,
        in1(1) => S1337,
        out1 => S1517
    );
notg_2090: ENTITY WORK.notg
    PORT MAP (
        in1 => S1517,
        out1 => S1518
    );
nor_n_2091: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1518,
        in1(1) => S1515,
        out1 => S1519
    );
nand_n_2092: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1517,
        in1(1) => S1516,
        out1 => S1520
    );
nand_n_2093: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1519,
        in1(1) => S202,
        out1 => S1521
    );
nand_n_2094: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1520,
        in1(1) => S203,
        out1 => S1522
    );
nor_n_2095: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1408,
        in1(1) => S1405,
        out1 => S1523
    );
nor_n_2096: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1523,
        in1(1) => S1410,
        out1 => S1524
    );
nor_n_2097: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1524,
        in1(1) => S1452,
        out1 => S1525
    );
nor_n_2098: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1453,
        in1(1) => S1350,
        out1 => S1526
    );
nor_n_2099: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1526,
        in1(1) => S1525,
        out1 => S1527
    );
notg_2100: ENTITY WORK.notg
    PORT MAP (
        in1 => S1527,
        out1 => S1528
    );
nor_n_2101: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1528,
        in1(1) => S209,
        out1 => S1529
    );
nand_n_2102: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1527,
        in1(1) => S208,
        out1 => S1530
    );
nor_n_2103: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1453,
        in1(1) => S1360,
        out1 => S1531
    );
nand_n_2104: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1452,
        in1(1) => S1361,
        out1 => S1532
    );
nor_n_2105: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1401,
        in1(1) => S1366,
        out1 => S1533
    );
nor_n_2106: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1533,
        in1(1) => S1402,
        out1 => S1534
    );
nor_n_2107: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1534,
        in1(1) => S1452,
        out1 => S1535
    );
notg_2108: ENTITY WORK.notg
    PORT MAP (
        in1 => S1535,
        out1 => S1536
    );
nor_n_2109: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1535,
        in1(1) => S1531,
        out1 => S1537
    );
nand_n_2110: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1536,
        in1(1) => S1532,
        out1 => S1538
    );
nor_n_2111: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1538,
        in1(1) => S241,
        out1 => S1539
    );
nand_n_2112: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1537,
        in1(1) => S240,
        out1 => S1540
    );
nor_n_2113: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1537,
        in1(1) => S240,
        out1 => S1541
    );
nand_n_2114: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1538,
        in1(1) => S241,
        out1 => S1542
    );
nor_n_2115: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1541,
        in1(1) => S1539,
        out1 => S1543
    );
nand_n_2116: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1542,
        in1(1) => S1540,
        out1 => S1544
    );
nand_n_2117: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1396,
        in1(1) => S1381,
        out1 => S1545
    );
nand_n_2118: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1545,
        in1(1) => S1399,
        out1 => S1546
    );
nand_n_2119: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1546,
        in1(1) => S1453,
        out1 => S1547
    );
nand_n_2120: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1452,
        in1(1) => S1375,
        out1 => S1548
    );
nand_n_2121: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1548,
        in1(1) => S1547,
        out1 => S1549
    );
notg_2122: ENTITY WORK.notg
    PORT MAP (
        in1 => S1549,
        out1 => S1550
    );
nor_n_2123: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1549,
        in1(1) => S249,
        out1 => S1551
    );
nand_n_2124: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1550,
        in1(1) => S248,
        out1 => S1552
    );
nand_n_2125: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1549,
        in1(1) => S249,
        out1 => S1553
    );
nand_n_2126: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1553,
        in1(1) => S1552,
        out1 => S1554
    );
notg_2127: ENTITY WORK.notg
    PORT MAP (
        in1 => S1554,
        out1 => S1555
    );
nor_n_2128: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1392,
        in1(1) => S1203,
        out1 => S1556
    );
nor_n_2129: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1556,
        in1(1) => S1394,
        out1 => S1557
    );
nor_n_2130: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1557,
        in1(1) => S1452,
        out1 => S1558
    );
nor_n_2131: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1453,
        in1(1) => S1386,
        out1 => S1559
    );
nor_n_2132: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1559,
        in1(1) => S1558,
        out1 => S1560
    );
notg_2133: ENTITY WORK.notg
    PORT MAP (
        in1 => S1560,
        out1 => S1561
    );
nor_n_2134: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1561,
        in1(1) => S257,
        out1 => S1562
    );
nand_n_2135: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1560,
        in1(1) => S256,
        out1 => S1563
    );
nor_n_2136: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1560,
        in1(1) => S256,
        out1 => S1564
    );
nand_n_2137: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1561,
        in1(1) => S257,
        out1 => S1565
    );
nor_n_2138: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1452,
        in1(1) => S270,
        out1 => S1566
    );
nand_n_2139: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1453,
        in1(1) => S271,
        out1 => S1567
    );
nor_n_2140: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1566,
        in1(1) => S5936,
        out1 => S1568
    );
nand_n_2141: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1567,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S1569
    );
nor_n_2142: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1452,
        in1(1) => S1203,
        out1 => S1570
    );
nand_n_2143: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1453,
        in1(1) => S1202,
        out1 => S1571
    );
nor_n_2144: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1570,
        in1(1) => S1568,
        out1 => S1572
    );
nand_n_2145: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1571,
        in1(1) => S1569,
        out1 => S1573
    );
nor_n_2146: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1572,
        in1(1) => S265,
        out1 => S1574
    );
nand_n_2147: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1573,
        in1(1) => S264,
        out1 => S1575
    );
nor_n_2148: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1573,
        in1(1) => S264,
        out1 => S1576
    );
nand_n_2149: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1572,
        in1(1) => S265,
        out1 => S1577
    );
nor_n_2150: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1576,
        in1(1) => S1574,
        out1 => S1578
    );
nand_n_2151: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1577,
        in1(1) => S1575,
        out1 => S1579
    );
nor_n_2152: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S1580
    );
nand_n_2153: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => S5947,
        out1 => S1581
    );
nor_n_2154: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1580,
        in1(1) => S1579,
        out1 => S1582
    );
nand_n_2155: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1581,
        in1(1) => S1578,
        out1 => S1583
    );
nor_n_2156: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1582,
        in1(1) => S1574,
        out1 => S1584
    );
nand_n_2157: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1583,
        in1(1) => S1575,
        out1 => S1585
    );
nor_n_2158: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1584,
        in1(1) => S1564,
        out1 => S1586
    );
nand_n_2159: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1585,
        in1(1) => S1565,
        out1 => S1587
    );
nor_n_2160: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1586,
        in1(1) => S1562,
        out1 => S1588
    );
nand_n_2161: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1587,
        in1(1) => S1563,
        out1 => S1589
    );
nor_n_2162: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1588,
        in1(1) => S1554,
        out1 => S1590
    );
nand_n_2163: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1589,
        in1(1) => S1555,
        out1 => S1591
    );
nor_n_2164: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1590,
        in1(1) => S1551,
        out1 => S1592
    );
nand_n_2165: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1591,
        in1(1) => S1552,
        out1 => S1593
    );
nor_n_2166: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1592,
        in1(1) => S1544,
        out1 => S1594
    );
nand_n_2167: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1593,
        in1(1) => S1543,
        out1 => S1595
    );
nor_n_2168: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1594,
        in1(1) => S1539,
        out1 => S1596
    );
nand_n_2169: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1595,
        in1(1) => S1540,
        out1 => S1597
    );
nor_n_2170: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1527,
        in1(1) => S208,
        out1 => S1598
    );
nor_n_2171: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1598,
        in1(1) => S1529,
        out1 => S1599
    );
notg_2172: ENTITY WORK.notg
    PORT MAP (
        in1 => S1599,
        out1 => S1600
    );
nor_n_2173: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1600,
        in1(1) => S1596,
        out1 => S1601
    );
nand_n_2174: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1599,
        in1(1) => S1597,
        out1 => S1602
    );
nor_n_2175: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1601,
        in1(1) => S1529,
        out1 => S1603
    );
nand_n_2176: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1602,
        in1(1) => S1530,
        out1 => S1604
    );
nand_n_2177: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1604,
        in1(1) => S1522,
        out1 => S1605
    );
nand_n_2178: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1603,
        in1(1) => S1521,
        out1 => S1606
    );
nand_n_2179: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1606,
        in1(1) => S1522,
        out1 => S1607
    );
nand_n_2180: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1605,
        in1(1) => S1521,
        out1 => S1608
    );
nor_n_2181: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1607,
        in1(1) => S1511,
        out1 => S1609
    );
nand_n_2182: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1608,
        in1(1) => S1512,
        out1 => S1610
    );
nor_n_2183: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1609,
        in1(1) => S1508,
        out1 => S1611
    );
nand_n_2184: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1610,
        in1(1) => S1509,
        out1 => S1612
    );
nor_n_2185: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1611,
        in1(1) => S1501,
        out1 => S1613
    );
nor_n_2186: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1612,
        in1(1) => S1500,
        out1 => S1614
    );
nor_n_2187: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1613,
        in1(1) => S1500,
        out1 => S1615
    );
nor_n_2188: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1614,
        in1(1) => S1501,
        out1 => S1616
    );
nor_n_2189: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1615,
        in1(1) => S1487,
        out1 => S1617
    );
nand_n_2190: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1616,
        in1(1) => S1488,
        out1 => S1618
    );
nor_n_2191: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1617,
        in1(1) => S1484,
        out1 => S1619
    );
nand_n_2192: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1618,
        in1(1) => S1485,
        out1 => S1620
    );
nor_n_2193: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1620,
        in1(1) => S1477,
        out1 => S1621
    );
nor_n_2194: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1619,
        in1(1) => S1476,
        out1 => S1622
    );
nor_n_2195: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1621,
        in1(1) => S1476,
        out1 => S1623
    );
nor_n_2196: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1622,
        in1(1) => S1477,
        out1 => S1624
    );
nor_n_2197: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1624,
        in1(1) => S1463,
        out1 => S1625
    );
nand_n_2198: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1623,
        in1(1) => S1464,
        out1 => S1626
    );
nor_n_2199: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1625,
        in1(1) => S1460,
        out1 => S1627
    );
nand_n_2200: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1626,
        in1(1) => S1461,
        out1 => S1628
    );
nor_n_2201: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1628,
        in1(1) => S1443,
        out1 => S1629
    );
nand_n_2202: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1627,
        in1(1) => S1444,
        out1 => S1630
    );
nand_n_2203: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1258,
        in1(1) => new_datapath_multdivunit_1697_B_12,
        out1 => S1631
    );
nand_n_2204: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1631,
        in1(1) => S212,
        out1 => S1632
    );
notg_2205: ENTITY WORK.notg
    PORT MAP (
        in1 => S1632,
        out1 => S1633
    );
nor_n_2206: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1632,
        in1(1) => S1629,
        out1 => S1634
    );
nand_n_2207: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1633,
        in1(1) => S1630,
        out1 => S1635
    );
nand_n_2208: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1624,
        in1(1) => S1463,
        out1 => S1636
    );
nand_n_2209: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1636,
        in1(1) => S1626,
        out1 => S1637
    );
nand_n_2210: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1637,
        in1(1) => S1634,
        out1 => S1638
    );
nand_n_2211: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1635,
        in1(1) => S1458,
        out1 => S1639
    );
nand_n_2212: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1639,
        in1(1) => S1638,
        out1 => S1640
    );
notg_2213: ENTITY WORK.notg
    PORT MAP (
        in1 => S1640,
        out1 => S1641
    );
nor_n_2214: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1640,
        in1(1) => new_datapath_multdivunit_1697_B_12,
        out1 => S1642
    );
nand_n_2215: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1641,
        in1(1) => S3434,
        out1 => S1643
    );
nand_n_2216: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1640,
        in1(1) => new_datapath_multdivunit_1697_B_12,
        out1 => S1644
    );
nand_n_2217: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1644,
        in1(1) => S1643,
        out1 => S1645
    );
notg_2218: ENTITY WORK.notg
    PORT MAP (
        in1 => S1645,
        out1 => S1646
    );
nor_n_2219: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1477,
        in1(1) => S1476,
        out1 => S1647
    );
nor_n_2220: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1647,
        in1(1) => S1620,
        out1 => S1648
    );
notg_2221: ENTITY WORK.notg
    PORT MAP (
        in1 => S1648,
        out1 => S1649
    );
nand_n_2222: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1647,
        in1(1) => S1620,
        out1 => S1650
    );
notg_2223: ENTITY WORK.notg
    PORT MAP (
        in1 => S1650,
        out1 => S1651
    );
nor_n_2224: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1651,
        in1(1) => S1648,
        out1 => S1652
    );
nand_n_2225: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1650,
        in1(1) => S1649,
        out1 => S1653
    );
nor_n_2226: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1652,
        in1(1) => S1635,
        out1 => S1654
    );
nand_n_2227: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1653,
        in1(1) => S1634,
        out1 => S1655
    );
nor_n_2228: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1634,
        in1(1) => S1475,
        out1 => S1656
    );
nand_n_2229: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1635,
        in1(1) => S1474,
        out1 => S1657
    );
nor_n_2230: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1656,
        in1(1) => S1654,
        out1 => S1658
    );
nand_n_2231: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1657,
        in1(1) => S1655,
        out1 => S1659
    );
nor_n_2232: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1659,
        in1(1) => new_datapath_multdivunit_1697_B_11,
        out1 => S1660
    );
nand_n_2233: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1658,
        in1(1) => S3445,
        out1 => S1661
    );
nor_n_2234: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1658,
        in1(1) => S3445,
        out1 => S1662
    );
nand_n_2235: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1659,
        in1(1) => new_datapath_multdivunit_1697_B_11,
        out1 => S1663
    );
nand_n_2236: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1615,
        in1(1) => S1487,
        out1 => S1664
    );
nand_n_2237: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1664,
        in1(1) => S1618,
        out1 => S1665
    );
nand_n_2238: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1665,
        in1(1) => S1634,
        out1 => S1666
    );
nand_n_2239: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1635,
        in1(1) => S1482,
        out1 => S1667
    );
nand_n_2240: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1667,
        in1(1) => S1666,
        out1 => S1668
    );
notg_2241: ENTITY WORK.notg
    PORT MAP (
        in1 => S1668,
        out1 => S1669
    );
nor_n_2242: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1668,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S1670
    );
nand_n_2243: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1669,
        in1(1) => S3456,
        out1 => S1671
    );
nand_n_2244: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1668,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S1672
    );
notg_2245: ENTITY WORK.notg
    PORT MAP (
        in1 => S1672,
        out1 => S1673
    );
nor_n_2246: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1673,
        in1(1) => S1670,
        out1 => S1674
    );
nand_n_2247: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1672,
        in1(1) => S1671,
        out1 => S1675
    );
nor_n_2248: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1501,
        in1(1) => S1500,
        out1 => S1676
    );
nor_n_2249: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1676,
        in1(1) => S1612,
        out1 => S1677
    );
notg_2250: ENTITY WORK.notg
    PORT MAP (
        in1 => S1677,
        out1 => S1678
    );
nand_n_2251: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1676,
        in1(1) => S1612,
        out1 => S1679
    );
notg_2252: ENTITY WORK.notg
    PORT MAP (
        in1 => S1679,
        out1 => S1680
    );
nor_n_2253: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1680,
        in1(1) => S1677,
        out1 => S1681
    );
nand_n_2254: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1679,
        in1(1) => S1678,
        out1 => S1682
    );
nor_n_2255: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1681,
        in1(1) => S1635,
        out1 => S1683
    );
nand_n_2256: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1682,
        in1(1) => S1634,
        out1 => S1684
    );
nor_n_2257: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1634,
        in1(1) => S1498,
        out1 => S1685
    );
nand_n_2258: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1635,
        in1(1) => S1499,
        out1 => S1686
    );
nor_n_2259: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1685,
        in1(1) => S1683,
        out1 => S1687
    );
nand_n_2260: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1686,
        in1(1) => S1684,
        out1 => S1688
    );
nand_n_2261: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1687,
        in1(1) => S3467,
        out1 => S1689
    );
nand_n_2262: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1688,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S1690
    );
nand_n_2263: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1607,
        in1(1) => S1511,
        out1 => S1691
    );
nand_n_2264: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1691,
        in1(1) => S1610,
        out1 => S1692
    );
nand_n_2265: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1692,
        in1(1) => S1634,
        out1 => S1693
    );
nand_n_2266: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1635,
        in1(1) => S1506,
        out1 => S1694
    );
nand_n_2267: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1694,
        in1(1) => S1693,
        out1 => S1695
    );
notg_2268: ENTITY WORK.notg
    PORT MAP (
        in1 => S1695,
        out1 => S1696
    );
nor_n_2269: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1695,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S1697
    );
nand_n_2270: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1696,
        in1(1) => S3478,
        out1 => S1698
    );
nand_n_2271: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1695,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S1699
    );
nand_n_2272: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1699,
        in1(1) => S1698,
        out1 => S1700
    );
notg_2273: ENTITY WORK.notg
    PORT MAP (
        in1 => S1700,
        out1 => S1701
    );
nand_n_2274: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1522,
        in1(1) => S1521,
        out1 => S1702
    );
nand_n_2275: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1702,
        in1(1) => S1603,
        out1 => S1703
    );
notg_2276: ENTITY WORK.notg
    PORT MAP (
        in1 => S1703,
        out1 => S1704
    );
nor_n_2277: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1702,
        in1(1) => S1603,
        out1 => S1705
    );
nor_n_2278: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1705,
        in1(1) => S1704,
        out1 => S1706
    );
nor_n_2279: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1706,
        in1(1) => S1635,
        out1 => S1707
    );
nor_n_2280: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1634,
        in1(1) => S1519,
        out1 => S1708
    );
nor_n_2281: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1708,
        in1(1) => S1707,
        out1 => S1709
    );
notg_2282: ENTITY WORK.notg
    PORT MAP (
        in1 => S1709,
        out1 => S1710
    );
nand_n_2283: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1709,
        in1(1) => S228,
        out1 => S1711
    );
nand_n_2284: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1710,
        in1(1) => S229,
        out1 => S1712
    );
nor_n_2285: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1599,
        in1(1) => S1597,
        out1 => S1713
    );
nor_n_2286: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1713,
        in1(1) => S1601,
        out1 => S1714
    );
nor_n_2287: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1714,
        in1(1) => S1635,
        out1 => S1715
    );
nor_n_2288: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1634,
        in1(1) => S1527,
        out1 => S1716
    );
nor_n_2289: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1716,
        in1(1) => S1715,
        out1 => S1717
    );
notg_2290: ENTITY WORK.notg
    PORT MAP (
        in1 => S1717,
        out1 => S1718
    );
nor_n_2291: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1718,
        in1(1) => S203,
        out1 => S1719
    );
notg_2292: ENTITY WORK.notg
    PORT MAP (
        in1 => S1719,
        out1 => S1720
    );
nor_n_2293: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1593,
        in1(1) => S1543,
        out1 => S1721
    );
notg_2294: ENTITY WORK.notg
    PORT MAP (
        in1 => S1721,
        out1 => S1722
    );
nor_n_2295: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1721,
        in1(1) => S1594,
        out1 => S1723
    );
nand_n_2296: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1722,
        in1(1) => S1595,
        out1 => S1724
    );
nor_n_2297: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1723,
        in1(1) => S1635,
        out1 => S1725
    );
nand_n_2298: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1724,
        in1(1) => S1634,
        out1 => S1726
    );
nor_n_2299: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1634,
        in1(1) => S1537,
        out1 => S1727
    );
nand_n_2300: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1635,
        in1(1) => S1538,
        out1 => S1728
    );
nor_n_2301: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1727,
        in1(1) => S1725,
        out1 => S1729
    );
nand_n_2302: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1728,
        in1(1) => S1726,
        out1 => S1730
    );
nor_n_2303: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1730,
        in1(1) => S209,
        out1 => S1731
    );
nand_n_2304: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1729,
        in1(1) => S208,
        out1 => S1732
    );
nor_n_2305: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1729,
        in1(1) => S208,
        out1 => S1733
    );
nor_n_2306: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1733,
        in1(1) => S1731,
        out1 => S1734
    );
notg_2307: ENTITY WORK.notg
    PORT MAP (
        in1 => S1734,
        out1 => S1735
    );
nand_n_2308: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1588,
        in1(1) => S1554,
        out1 => S1736
    );
nand_n_2309: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1736,
        in1(1) => S1591,
        out1 => S1737
    );
nand_n_2310: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1737,
        in1(1) => S1634,
        out1 => S1738
    );
nand_n_2311: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1635,
        in1(1) => S1549,
        out1 => S1739
    );
nand_n_2312: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1739,
        in1(1) => S1738,
        out1 => S1740
    );
notg_2313: ENTITY WORK.notg
    PORT MAP (
        in1 => S1740,
        out1 => S1741
    );
nand_n_2314: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1741,
        in1(1) => S240,
        out1 => S1742
    );
notg_2315: ENTITY WORK.notg
    PORT MAP (
        in1 => S1742,
        out1 => S1743
    );
nand_n_2316: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1740,
        in1(1) => S241,
        out1 => S1744
    );
nand_n_2317: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1744,
        in1(1) => S1742,
        out1 => S1745
    );
notg_2318: ENTITY WORK.notg
    PORT MAP (
        in1 => S1745,
        out1 => S1746
    );
nor_n_2319: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1564,
        in1(1) => S1562,
        out1 => S1747
    );
nand_n_2320: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1565,
        in1(1) => S1563,
        out1 => S1748
    );
nand_n_2321: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1747,
        in1(1) => S1584,
        out1 => S1749
    );
nand_n_2322: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1748,
        in1(1) => S1585,
        out1 => S1750
    );
nand_n_2323: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1750,
        in1(1) => S1749,
        out1 => S1751
    );
nand_n_2324: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1751,
        in1(1) => S1634,
        out1 => S1752
    );
nand_n_2325: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1635,
        in1(1) => S1560,
        out1 => S1753
    );
nand_n_2326: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1753,
        in1(1) => S1752,
        out1 => S1754
    );
notg_2327: ENTITY WORK.notg
    PORT MAP (
        in1 => S1754,
        out1 => S1755
    );
nor_n_2328: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1755,
        in1(1) => S249,
        out1 => S1756
    );
notg_2329: ENTITY WORK.notg
    PORT MAP (
        in1 => S1756,
        out1 => S1757
    );
nor_n_2330: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1754,
        in1(1) => S248,
        out1 => S1758
    );
nor_n_2331: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1758,
        in1(1) => S1756,
        out1 => S1759
    );
notg_2332: ENTITY WORK.notg
    PORT MAP (
        in1 => S1759,
        out1 => S1760
    );
nor_n_2333: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1581,
        in1(1) => S1578,
        out1 => S1761
    );
nand_n_2334: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1580,
        in1(1) => S1579,
        out1 => S1762
    );
nor_n_2335: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1761,
        in1(1) => S1582,
        out1 => S1763
    );
nand_n_2336: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1762,
        in1(1) => S1583,
        out1 => S1764
    );
nor_n_2337: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1763,
        in1(1) => S1635,
        out1 => S1765
    );
nand_n_2338: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1764,
        in1(1) => S1634,
        out1 => S1766
    );
nor_n_2339: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1634,
        in1(1) => S1573,
        out1 => S1767
    );
nand_n_2340: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1635,
        in1(1) => S1572,
        out1 => S1768
    );
nor_n_2341: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1767,
        in1(1) => S1765,
        out1 => S1769
    );
nand_n_2342: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1768,
        in1(1) => S1766,
        out1 => S1770
    );
nor_n_2343: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1770,
        in1(1) => S257,
        out1 => S1771
    );
nand_n_2344: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1769,
        in1(1) => S256,
        out1 => S1772
    );
nor_n_2345: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1769,
        in1(1) => S256,
        out1 => S1773
    );
nand_n_2346: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1770,
        in1(1) => S257,
        out1 => S1774
    );
nor_n_2347: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1773,
        in1(1) => S1771,
        out1 => S1775
    );
nand_n_2348: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1774,
        in1(1) => S1772,
        out1 => S1776
    );
nor_n_2349: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1635,
        in1(1) => S270,
        out1 => S1777
    );
nand_n_2350: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1634,
        in1(1) => S271,
        out1 => S1778
    );
nor_n_2351: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1777,
        in1(1) => S5947,
        out1 => S1779
    );
nand_n_2352: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1778,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S1780
    );
nor_n_2353: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1635,
        in1(1) => S1581,
        out1 => S1781
    );
nand_n_2354: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1634,
        in1(1) => S1580,
        out1 => S1782
    );
nor_n_2355: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1781,
        in1(1) => S1779,
        out1 => S1783
    );
nand_n_2356: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1782,
        in1(1) => S1780,
        out1 => S1784
    );
nor_n_2357: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1783,
        in1(1) => S265,
        out1 => S1785
    );
nand_n_2358: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1784,
        in1(1) => S264,
        out1 => S1786
    );
nor_n_2359: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S1787
    );
nand_n_2360: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => S5957,
        out1 => S1788
    );
nor_n_2361: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1784,
        in1(1) => S264,
        out1 => S1789
    );
nand_n_2362: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1783,
        in1(1) => S265,
        out1 => S1790
    );
nor_n_2363: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1789,
        in1(1) => S1785,
        out1 => S1791
    );
nand_n_2364: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1790,
        in1(1) => S1786,
        out1 => S1792
    );
nor_n_2365: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1792,
        in1(1) => S1787,
        out1 => S1793
    );
nand_n_2366: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1791,
        in1(1) => S1788,
        out1 => S1794
    );
nor_n_2367: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1793,
        in1(1) => S1785,
        out1 => S1795
    );
nand_n_2368: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1794,
        in1(1) => S1786,
        out1 => S1796
    );
nor_n_2369: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1795,
        in1(1) => S1776,
        out1 => S1797
    );
nand_n_2370: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1796,
        in1(1) => S1775,
        out1 => S1798
    );
nor_n_2371: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1797,
        in1(1) => S1771,
        out1 => S1799
    );
nand_n_2372: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1798,
        in1(1) => S1772,
        out1 => S1800
    );
nor_n_2373: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1799,
        in1(1) => S1760,
        out1 => S1801
    );
nand_n_2374: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1800,
        in1(1) => S1759,
        out1 => S1802
    );
nor_n_2375: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1801,
        in1(1) => S1756,
        out1 => S1803
    );
nand_n_2376: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1802,
        in1(1) => S1757,
        out1 => S1804
    );
nor_n_2377: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1803,
        in1(1) => S1745,
        out1 => S1805
    );
nand_n_2378: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1804,
        in1(1) => S1746,
        out1 => S1806
    );
nor_n_2379: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1805,
        in1(1) => S1743,
        out1 => S1807
    );
nand_n_2380: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1806,
        in1(1) => S1742,
        out1 => S1808
    );
nor_n_2381: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1807,
        in1(1) => S1735,
        out1 => S1809
    );
nand_n_2382: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1808,
        in1(1) => S1734,
        out1 => S1810
    );
nor_n_2383: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1809,
        in1(1) => S1731,
        out1 => S1811
    );
nand_n_2384: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1810,
        in1(1) => S1732,
        out1 => S1812
    );
nor_n_2385: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1717,
        in1(1) => S202,
        out1 => S1813
    );
nor_n_2386: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1813,
        in1(1) => S1719,
        out1 => S1814
    );
notg_2387: ENTITY WORK.notg
    PORT MAP (
        in1 => S1814,
        out1 => S1815
    );
nor_n_2388: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1815,
        in1(1) => S1811,
        out1 => S1816
    );
nand_n_2389: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1814,
        in1(1) => S1812,
        out1 => S1817
    );
nor_n_2390: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1816,
        in1(1) => S1719,
        out1 => S1818
    );
nand_n_2391: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1817,
        in1(1) => S1720,
        out1 => S1819
    );
nand_n_2392: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1819,
        in1(1) => S1712,
        out1 => S1820
    );
nand_n_2393: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1818,
        in1(1) => S1711,
        out1 => S1821
    );
nand_n_2394: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1821,
        in1(1) => S1712,
        out1 => S1822
    );
nand_n_2395: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1820,
        in1(1) => S1711,
        out1 => S1823
    );
nor_n_2396: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1822,
        in1(1) => S1700,
        out1 => S1824
    );
nand_n_2397: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1823,
        in1(1) => S1701,
        out1 => S1825
    );
nor_n_2398: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1824,
        in1(1) => S1697,
        out1 => S1826
    );
nand_n_2399: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1825,
        in1(1) => S1698,
        out1 => S1827
    );
nand_n_2400: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1827,
        in1(1) => S1690,
        out1 => S1828
    );
nand_n_2401: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1826,
        in1(1) => S1689,
        out1 => S1829
    );
nand_n_2402: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1829,
        in1(1) => S1690,
        out1 => S1830
    );
nand_n_2403: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1828,
        in1(1) => S1689,
        out1 => S1831
    );
nor_n_2404: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1830,
        in1(1) => S1675,
        out1 => S1832
    );
nand_n_2405: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1831,
        in1(1) => S1674,
        out1 => S1833
    );
nor_n_2406: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1832,
        in1(1) => S1670,
        out1 => S1834
    );
nand_n_2407: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1833,
        in1(1) => S1671,
        out1 => S1835
    );
nor_n_2408: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1834,
        in1(1) => S1662,
        out1 => S1836
    );
nand_n_2409: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1835,
        in1(1) => S1663,
        out1 => S1837
    );
nor_n_2410: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1836,
        in1(1) => S1660,
        out1 => S1838
    );
nand_n_2411: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1837,
        in1(1) => S1661,
        out1 => S1839
    );
nor_n_2412: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1838,
        in1(1) => S1645,
        out1 => S1840
    );
nand_n_2413: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1839,
        in1(1) => S1646,
        out1 => S1841
    );
nor_n_2414: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1840,
        in1(1) => S1642,
        out1 => S1842
    );
nand_n_2415: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1841,
        in1(1) => S1643,
        out1 => S1843
    );
nand_n_2416: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S212,
        in1(1) => new_datapath_multdivunit_1697_B_12,
        out1 => S1844
    );
nand_n_2417: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1627,
        in1(1) => S214,
        out1 => S1845
    );
nor_n_2418: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1844,
        in1(1) => S1627,
        out1 => S1846
    );
nor_n_2419: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1846,
        in1(1) => S1442,
        out1 => S1847
    );
nand_n_2420: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1847,
        in1(1) => S1845,
        out1 => S1848
    );
nor_n_2421: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1848,
        in1(1) => new_datapath_multdivunit_1697_B_13,
        out1 => S1849
    );
notg_2422: ENTITY WORK.notg
    PORT MAP (
        in1 => S1849,
        out1 => S1850
    );
nor_n_2423: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1849,
        in1(1) => S1843,
        out1 => S1851
    );
nand_n_2424: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1850,
        in1(1) => S1842,
        out1 => S1852
    );
nand_n_2425: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1442,
        in1(1) => new_datapath_multdivunit_1697_B_13,
        out1 => S1853
    );
nand_n_2426: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1853,
        in1(1) => S210,
        out1 => S1854
    );
notg_2427: ENTITY WORK.notg
    PORT MAP (
        in1 => S1854,
        out1 => S1855
    );
nor_n_2428: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1854,
        in1(1) => S1851,
        out1 => S1856
    );
nand_n_2429: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1855,
        in1(1) => S1852,
        out1 => S1857
    );
nand_n_2430: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1838,
        in1(1) => S1645,
        out1 => S1858
    );
nand_n_2431: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1858,
        in1(1) => S1841,
        out1 => S1859
    );
nand_n_2432: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1859,
        in1(1) => S1856,
        out1 => S1860
    );
nand_n_2433: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1857,
        in1(1) => S1640,
        out1 => S1861
    );
nand_n_2434: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1861,
        in1(1) => S1860,
        out1 => S1862
    );
notg_2435: ENTITY WORK.notg
    PORT MAP (
        in1 => S1862,
        out1 => S1863
    );
nor_n_2436: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1862,
        in1(1) => new_datapath_multdivunit_1697_B_13,
        out1 => S1864
    );
nand_n_2437: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1863,
        in1(1) => S3423,
        out1 => S1865
    );
nand_n_2438: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1862,
        in1(1) => new_datapath_multdivunit_1697_B_13,
        out1 => S1866
    );
nand_n_2439: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1866,
        in1(1) => S1865,
        out1 => S1867
    );
notg_2440: ENTITY WORK.notg
    PORT MAP (
        in1 => S1867,
        out1 => S1868
    );
nor_n_2441: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1662,
        in1(1) => S1660,
        out1 => S1869
    );
nand_n_2442: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1663,
        in1(1) => S1661,
        out1 => S1870
    );
nor_n_2443: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1869,
        in1(1) => S1835,
        out1 => S1871
    );
nor_n_2444: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1870,
        in1(1) => S1834,
        out1 => S1872
    );
nor_n_2445: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1872,
        in1(1) => S1871,
        out1 => S1873
    );
nor_n_2446: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1873,
        in1(1) => S1857,
        out1 => S1874
    );
notg_2447: ENTITY WORK.notg
    PORT MAP (
        in1 => S1874,
        out1 => S1875
    );
nand_n_2448: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1857,
        in1(1) => S1659,
        out1 => S1876
    );
notg_2449: ENTITY WORK.notg
    PORT MAP (
        in1 => S1876,
        out1 => S1877
    );
nor_n_2450: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1877,
        in1(1) => S1874,
        out1 => S1878
    );
nand_n_2451: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1876,
        in1(1) => S1875,
        out1 => S1879
    );
nand_n_2452: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1878,
        in1(1) => S3434,
        out1 => S1880
    );
nand_n_2453: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1879,
        in1(1) => new_datapath_multdivunit_1697_B_12,
        out1 => S1881
    );
nand_n_2454: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1830,
        in1(1) => S1675,
        out1 => S1882
    );
notg_2455: ENTITY WORK.notg
    PORT MAP (
        in1 => S1882,
        out1 => S1883
    );
nor_n_2456: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1883,
        in1(1) => S1832,
        out1 => S1884
    );
nor_n_2457: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1884,
        in1(1) => S1857,
        out1 => S1885
    );
notg_2458: ENTITY WORK.notg
    PORT MAP (
        in1 => S1885,
        out1 => S1886
    );
nand_n_2459: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1857,
        in1(1) => S1668,
        out1 => S1887
    );
notg_2460: ENTITY WORK.notg
    PORT MAP (
        in1 => S1887,
        out1 => S1888
    );
nor_n_2461: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1888,
        in1(1) => S1885,
        out1 => S1889
    );
nand_n_2462: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1887,
        in1(1) => S1886,
        out1 => S1890
    );
nor_n_2463: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1890,
        in1(1) => new_datapath_multdivunit_1697_B_11,
        out1 => S1891
    );
notg_2464: ENTITY WORK.notg
    PORT MAP (
        in1 => S1891,
        out1 => S1892
    );
nand_n_2465: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1890,
        in1(1) => new_datapath_multdivunit_1697_B_11,
        out1 => S1893
    );
notg_2466: ENTITY WORK.notg
    PORT MAP (
        in1 => S1893,
        out1 => S1894
    );
nor_n_2467: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1894,
        in1(1) => S1891,
        out1 => S1895
    );
notg_2468: ENTITY WORK.notg
    PORT MAP (
        in1 => S1895,
        out1 => S1896
    );
nand_n_2469: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1690,
        in1(1) => S1689,
        out1 => S1897
    );
nand_n_2470: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1897,
        in1(1) => S1826,
        out1 => S1898
    );
notg_2471: ENTITY WORK.notg
    PORT MAP (
        in1 => S1898,
        out1 => S1899
    );
nor_n_2472: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1897,
        in1(1) => S1826,
        out1 => S1900
    );
nor_n_2473: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1900,
        in1(1) => S1899,
        out1 => S1901
    );
nor_n_2474: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1901,
        in1(1) => S1857,
        out1 => S1902
    );
notg_2475: ENTITY WORK.notg
    PORT MAP (
        in1 => S1902,
        out1 => S1903
    );
nand_n_2476: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1857,
        in1(1) => S1688,
        out1 => S1904
    );
notg_2477: ENTITY WORK.notg
    PORT MAP (
        in1 => S1904,
        out1 => S1905
    );
nor_n_2478: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1905,
        in1(1) => S1902,
        out1 => S1906
    );
nand_n_2479: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1904,
        in1(1) => S1903,
        out1 => S1907
    );
nand_n_2480: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1906,
        in1(1) => S3456,
        out1 => S1908
    );
nand_n_2481: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1907,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S1909
    );
nand_n_2482: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1822,
        in1(1) => S1700,
        out1 => S1910
    );
nand_n_2483: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1910,
        in1(1) => S1825,
        out1 => S1911
    );
nand_n_2484: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1911,
        in1(1) => S1856,
        out1 => S1912
    );
nand_n_2485: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1857,
        in1(1) => S1695,
        out1 => S1913
    );
nand_n_2486: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1913,
        in1(1) => S1912,
        out1 => S1914
    );
notg_2487: ENTITY WORK.notg
    PORT MAP (
        in1 => S1914,
        out1 => S1915
    );
nor_n_2488: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1914,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S1916
    );
nand_n_2489: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1915,
        in1(1) => S3467,
        out1 => S1917
    );
nand_n_2490: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1914,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S1918
    );
nand_n_2491: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1918,
        in1(1) => S1917,
        out1 => S1919
    );
notg_2492: ENTITY WORK.notg
    PORT MAP (
        in1 => S1919,
        out1 => S1920
    );
nand_n_2493: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1712,
        in1(1) => S1711,
        out1 => S1921
    );
nand_n_2494: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1921,
        in1(1) => S1818,
        out1 => S1922
    );
notg_2495: ENTITY WORK.notg
    PORT MAP (
        in1 => S1922,
        out1 => S1923
    );
nor_n_2496: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1921,
        in1(1) => S1818,
        out1 => S1924
    );
nor_n_2497: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1924,
        in1(1) => S1923,
        out1 => S1925
    );
nor_n_2498: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1925,
        in1(1) => S1857,
        out1 => S1926
    );
nand_n_2499: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1857,
        in1(1) => S1710,
        out1 => S1927
    );
notg_2500: ENTITY WORK.notg
    PORT MAP (
        in1 => S1927,
        out1 => S1928
    );
nor_n_2501: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1928,
        in1(1) => S1926,
        out1 => S1929
    );
notg_2502: ENTITY WORK.notg
    PORT MAP (
        in1 => S1929,
        out1 => S1930
    );
nand_n_2503: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1929,
        in1(1) => S3478,
        out1 => S1931
    );
nand_n_2504: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1930,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S1932
    );
nor_n_2505: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1814,
        in1(1) => S1812,
        out1 => S1933
    );
nor_n_2506: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1933,
        in1(1) => S1816,
        out1 => S1934
    );
nor_n_2507: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1934,
        in1(1) => S1857,
        out1 => S1935
    );
nor_n_2508: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1856,
        in1(1) => S1717,
        out1 => S1936
    );
nor_n_2509: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1936,
        in1(1) => S1935,
        out1 => S1937
    );
notg_2510: ENTITY WORK.notg
    PORT MAP (
        in1 => S1937,
        out1 => S1938
    );
nor_n_2511: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1938,
        in1(1) => S229,
        out1 => S1939
    );
notg_2512: ENTITY WORK.notg
    PORT MAP (
        in1 => S1939,
        out1 => S1940
    );
nor_n_2513: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1937,
        in1(1) => S228,
        out1 => S1941
    );
nor_n_2514: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1941,
        in1(1) => S1939,
        out1 => S1942
    );
notg_2515: ENTITY WORK.notg
    PORT MAP (
        in1 => S1942,
        out1 => S1943
    );
nand_n_2516: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1857,
        in1(1) => S1730,
        out1 => S1944
    );
notg_2517: ENTITY WORK.notg
    PORT MAP (
        in1 => S1944,
        out1 => S1945
    );
nor_n_2518: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1808,
        in1(1) => S1734,
        out1 => S1946
    );
nor_n_2519: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1946,
        in1(1) => S1809,
        out1 => S1947
    );
nor_n_2520: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1947,
        in1(1) => S1857,
        out1 => S1948
    );
notg_2521: ENTITY WORK.notg
    PORT MAP (
        in1 => S1948,
        out1 => S1949
    );
nor_n_2522: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1948,
        in1(1) => S1945,
        out1 => S1950
    );
nand_n_2523: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1949,
        in1(1) => S1944,
        out1 => S1951
    );
nor_n_2524: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1951,
        in1(1) => S203,
        out1 => S1952
    );
nor_n_2525: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1950,
        in1(1) => S202,
        out1 => S1953
    );
nand_n_2526: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1803,
        in1(1) => S1745,
        out1 => S1954
    );
nand_n_2527: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1954,
        in1(1) => S1806,
        out1 => S1955
    );
nand_n_2528: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1955,
        in1(1) => S1856,
        out1 => S1956
    );
nand_n_2529: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1857,
        in1(1) => S1740,
        out1 => S1957
    );
nand_n_2530: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1957,
        in1(1) => S1956,
        out1 => S1958
    );
notg_2531: ENTITY WORK.notg
    PORT MAP (
        in1 => S1958,
        out1 => S1959
    );
nand_n_2532: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1959,
        in1(1) => S208,
        out1 => S1960
    );
notg_2533: ENTITY WORK.notg
    PORT MAP (
        in1 => S1960,
        out1 => S1961
    );
nand_n_2534: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1958,
        in1(1) => S209,
        out1 => S1962
    );
nand_n_2535: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1962,
        in1(1) => S1960,
        out1 => S1963
    );
notg_2536: ENTITY WORK.notg
    PORT MAP (
        in1 => S1963,
        out1 => S1964
    );
nor_n_2537: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1800,
        in1(1) => S1759,
        out1 => S1965
    );
nor_n_2538: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1965,
        in1(1) => S1801,
        out1 => S1966
    );
nor_n_2539: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1966,
        in1(1) => S1857,
        out1 => S1967
    );
nor_n_2540: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1856,
        in1(1) => S1754,
        out1 => S1968
    );
nor_n_2541: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1968,
        in1(1) => S1967,
        out1 => S1969
    );
notg_2542: ENTITY WORK.notg
    PORT MAP (
        in1 => S1969,
        out1 => S1970
    );
nor_n_2543: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1970,
        in1(1) => S241,
        out1 => S1971
    );
nand_n_2544: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1969,
        in1(1) => S240,
        out1 => S1972
    );
nor_n_2545: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1969,
        in1(1) => S240,
        out1 => S1973
    );
nand_n_2546: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1970,
        in1(1) => S241,
        out1 => S1974
    );
nor_n_2547: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1796,
        in1(1) => S1775,
        out1 => S1975
    );
nor_n_2548: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1975,
        in1(1) => S1797,
        out1 => S1976
    );
nor_n_2549: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1976,
        in1(1) => S1857,
        out1 => S1977
    );
notg_2550: ENTITY WORK.notg
    PORT MAP (
        in1 => S1977,
        out1 => S1978
    );
nor_n_2551: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1856,
        in1(1) => S1769,
        out1 => S1979
    );
nand_n_2552: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1857,
        in1(1) => S1770,
        out1 => S1980
    );
nor_n_2553: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1979,
        in1(1) => S1977,
        out1 => S1981
    );
nand_n_2554: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1980,
        in1(1) => S1978,
        out1 => S1982
    );
nor_n_2555: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1982,
        in1(1) => S249,
        out1 => S1983
    );
nand_n_2556: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1981,
        in1(1) => S248,
        out1 => S1984
    );
nor_n_2557: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1981,
        in1(1) => S248,
        out1 => S1985
    );
nand_n_2558: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1982,
        in1(1) => S249,
        out1 => S1986
    );
nor_n_2559: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1985,
        in1(1) => S1983,
        out1 => S1987
    );
nand_n_2560: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1986,
        in1(1) => S1984,
        out1 => S1988
    );
nor_n_2561: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1791,
        in1(1) => S1788,
        out1 => S1989
    );
nor_n_2562: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1989,
        in1(1) => S1793,
        out1 => S1990
    );
nor_n_2563: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1990,
        in1(1) => S1857,
        out1 => S1991
    );
notg_2564: ENTITY WORK.notg
    PORT MAP (
        in1 => S1991,
        out1 => S1992
    );
nor_n_2565: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1856,
        in1(1) => S1784,
        out1 => S1993
    );
nand_n_2566: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1857,
        in1(1) => S1783,
        out1 => S1994
    );
nor_n_2567: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1993,
        in1(1) => S1991,
        out1 => S1995
    );
nand_n_2568: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1994,
        in1(1) => S1992,
        out1 => S1996
    );
nor_n_2569: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1996,
        in1(1) => S257,
        out1 => S1997
    );
nand_n_2570: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1995,
        in1(1) => S256,
        out1 => S1998
    );
nor_n_2571: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1995,
        in1(1) => S256,
        out1 => S1999
    );
nand_n_2572: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1996,
        in1(1) => S257,
        out1 => S2000
    );
nor_n_2573: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1999,
        in1(1) => S1997,
        out1 => S2001
    );
nand_n_2574: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2000,
        in1(1) => S1998,
        out1 => S2002
    );
nor_n_2575: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1857,
        in1(1) => S270,
        out1 => S2003
    );
nand_n_2576: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1856,
        in1(1) => S271,
        out1 => S2004
    );
nor_n_2577: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2004,
        in1(1) => S5957,
        out1 => S2005
    );
nand_n_2578: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2003,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S2006
    );
nor_n_2579: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2003,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S2007
    );
nand_n_2580: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2004,
        in1(1) => S5957,
        out1 => S2008
    );
nand_n_2581: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2008,
        in1(1) => S2006,
        out1 => S2009
    );
nor_n_2582: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2007,
        in1(1) => S2005,
        out1 => S2010
    );
nor_n_2583: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2009,
        in1(1) => S265,
        out1 => S2011
    );
nand_n_2584: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2010,
        in1(1) => S264,
        out1 => S2012
    );
nor_n_2585: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2010,
        in1(1) => S264,
        out1 => S2013
    );
nand_n_2586: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2009,
        in1(1) => S265,
        out1 => S2014
    );
nor_n_2587: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2013,
        in1(1) => S2011,
        out1 => S2015
    );
nand_n_2588: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2014,
        in1(1) => S2012,
        out1 => S2016
    );
nand_n_2589: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => S5966,
        out1 => S2017
    );
notg_2590: ENTITY WORK.notg
    PORT MAP (
        in1 => S2017,
        out1 => S2018
    );
nor_n_2591: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2018,
        in1(1) => S2016,
        out1 => S2019
    );
nand_n_2592: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2017,
        in1(1) => S2015,
        out1 => S2020
    );
nor_n_2593: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2019,
        in1(1) => S2011,
        out1 => S2021
    );
nand_n_2594: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2020,
        in1(1) => S2012,
        out1 => S2022
    );
nor_n_2595: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2021,
        in1(1) => S2002,
        out1 => S2023
    );
nand_n_2596: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2022,
        in1(1) => S2001,
        out1 => S2024
    );
nor_n_2597: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2023,
        in1(1) => S1997,
        out1 => S2025
    );
nand_n_2598: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2024,
        in1(1) => S1998,
        out1 => S2026
    );
nor_n_2599: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2025,
        in1(1) => S1988,
        out1 => S2027
    );
nand_n_2600: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2026,
        in1(1) => S1987,
        out1 => S2028
    );
nor_n_2601: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2027,
        in1(1) => S1983,
        out1 => S2029
    );
nand_n_2602: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2028,
        in1(1) => S1984,
        out1 => S2030
    );
nor_n_2603: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2029,
        in1(1) => S1973,
        out1 => S2031
    );
nand_n_2604: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2030,
        in1(1) => S1974,
        out1 => S2032
    );
nor_n_2605: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2031,
        in1(1) => S1971,
        out1 => S2033
    );
nand_n_2606: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2032,
        in1(1) => S1972,
        out1 => S2034
    );
nor_n_2607: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2033,
        in1(1) => S1963,
        out1 => S2035
    );
nand_n_2608: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2034,
        in1(1) => S1964,
        out1 => S2036
    );
nor_n_2609: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2035,
        in1(1) => S1961,
        out1 => S2037
    );
nand_n_2610: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2036,
        in1(1) => S1960,
        out1 => S2038
    );
nor_n_2611: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2037,
        in1(1) => S1953,
        out1 => S2039
    );
nor_n_2612: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2038,
        in1(1) => S1952,
        out1 => S2040
    );
nor_n_2613: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2039,
        in1(1) => S1952,
        out1 => S2041
    );
nor_n_2614: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2040,
        in1(1) => S1953,
        out1 => S2042
    );
nor_n_2615: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2041,
        in1(1) => S1943,
        out1 => S2043
    );
nand_n_2616: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2042,
        in1(1) => S1942,
        out1 => S2044
    );
nor_n_2617: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2043,
        in1(1) => S1939,
        out1 => S2045
    );
nand_n_2618: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2044,
        in1(1) => S1940,
        out1 => S2046
    );
nand_n_2619: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2046,
        in1(1) => S1932,
        out1 => S2047
    );
nand_n_2620: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2045,
        in1(1) => S1931,
        out1 => S2048
    );
nand_n_2621: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2048,
        in1(1) => S1932,
        out1 => S2049
    );
nand_n_2622: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2047,
        in1(1) => S1931,
        out1 => S2050
    );
nor_n_2623: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2049,
        in1(1) => S1919,
        out1 => S2051
    );
nand_n_2624: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2050,
        in1(1) => S1920,
        out1 => S2052
    );
nor_n_2625: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2051,
        in1(1) => S1916,
        out1 => S2053
    );
nand_n_2626: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2052,
        in1(1) => S1917,
        out1 => S2054
    );
nand_n_2627: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2054,
        in1(1) => S1909,
        out1 => S2055
    );
nand_n_2628: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2053,
        in1(1) => S1908,
        out1 => S2056
    );
nand_n_2629: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2056,
        in1(1) => S1909,
        out1 => S2057
    );
nand_n_2630: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2055,
        in1(1) => S1908,
        out1 => S2058
    );
nor_n_2631: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2057,
        in1(1) => S1896,
        out1 => S2059
    );
nand_n_2632: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2058,
        in1(1) => S1895,
        out1 => S2060
    );
nor_n_2633: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2059,
        in1(1) => S1891,
        out1 => S2061
    );
nand_n_2634: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2060,
        in1(1) => S1892,
        out1 => S2062
    );
nand_n_2635: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2062,
        in1(1) => S1881,
        out1 => S2063
    );
nand_n_2636: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2061,
        in1(1) => S1880,
        out1 => S2064
    );
nand_n_2637: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2064,
        in1(1) => S1881,
        out1 => S2065
    );
nand_n_2638: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2063,
        in1(1) => S1880,
        out1 => S2066
    );
nor_n_2639: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2065,
        in1(1) => S1867,
        out1 => S2067
    );
nand_n_2640: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2066,
        in1(1) => S1868,
        out1 => S2068
    );
nor_n_2641: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2067,
        in1(1) => S1864,
        out1 => S2069
    );
nand_n_2642: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2068,
        in1(1) => S1865,
        out1 => S2070
    );
nand_n_2643: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S210,
        in1(1) => new_datapath_multdivunit_1697_B_13,
        out1 => S2071
    );
nor_n_2644: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2071,
        in1(1) => S1842,
        out1 => S2072
    );
nand_n_2645: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1842,
        in1(1) => S212,
        out1 => S2073
    );
nor_n_2646: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2072,
        in1(1) => S1848,
        out1 => S2074
    );
nand_n_2647: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2074,
        in1(1) => S2073,
        out1 => S2075
    );
nor_n_2648: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2075,
        in1(1) => new_datapath_multdivunit_1697_B_14,
        out1 => S2076
    );
notg_2649: ENTITY WORK.notg
    PORT MAP (
        in1 => S2076,
        out1 => S2077
    );
nor_n_2650: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2076,
        in1(1) => S2070,
        out1 => S2078
    );
nand_n_2651: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2077,
        in1(1) => S2069,
        out1 => S2079
    );
nor_n_2652: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2075,
        in1(1) => new_datapath_multdivunit_1697_B_15,
        out1 => S2080
    );
nor_n_2653: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2080,
        in1(1) => S210,
        out1 => S2081
    );
notg_2654: ENTITY WORK.notg
    PORT MAP (
        in1 => S2081,
        out1 => S2082
    );
nor_n_2655: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2081,
        in1(1) => S2078,
        out1 => S2083
    );
nand_n_2656: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2082,
        in1(1) => S2079,
        out1 => S2084
    );
nand_n_2657: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2033,
        in1(1) => S1963,
        out1 => S2085
    );
nand_n_2658: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2085,
        in1(1) => S2036,
        out1 => S2086
    );
nand_n_2659: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2086,
        in1(1) => S2083,
        out1 => S2087
    );
nand_n_2660: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2084,
        in1(1) => S1958,
        out1 => S2088
    );
nand_n_2661: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2088,
        in1(1) => S2087,
        out1 => S2089
    );
nand_n_2662: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2089,
        in1(1) => S203,
        out1 => S2090
    );
nor_n_2663: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1973,
        in1(1) => S1971,
        out1 => S2091
    );
nand_n_2664: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1974,
        in1(1) => S1972,
        out1 => S2092
    );
nand_n_2665: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2091,
        in1(1) => S2029,
        out1 => S2093
    );
nand_n_2666: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2092,
        in1(1) => S2030,
        out1 => S2094
    );
nand_n_2667: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2094,
        in1(1) => S2093,
        out1 => S2095
    );
nor_n_2668: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2095,
        in1(1) => S2084,
        out1 => S2096
    );
nor_n_2669: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2083,
        in1(1) => S1969,
        out1 => S2097
    );
nor_n_2670: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2097,
        in1(1) => S2096,
        out1 => S2098
    );
nand_n_2671: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2098,
        in1(1) => S208,
        out1 => S2099
    );
nor_n_2672: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2017,
        in1(1) => S2015,
        out1 => S2100
    );
nor_n_2673: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2100,
        in1(1) => S2019,
        out1 => S2101
    );
nor_n_2674: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2101,
        in1(1) => S2084,
        out1 => S2102
    );
nor_n_2675: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2083,
        in1(1) => S2010,
        out1 => S2103
    );
nor_n_2676: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2103,
        in1(1) => S2102,
        out1 => S2104
    );
nand_n_2677: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2104,
        in1(1) => S256,
        out1 => S2105
    );
nand_n_2678: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2083,
        in1(1) => S271,
        out1 => S2106
    );
nand_n_2679: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2106,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S2107
    );
nor_n_2680: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S2108
    );
nor_n_2681: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2108,
        in1(1) => S265,
        out1 => S2109
    );
nor_n_2682: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2084,
        in1(1) => S2017,
        out1 => S2110
    );
nor_n_2683: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2110,
        in1(1) => S2109,
        out1 => S2111
    );
nand_n_2684: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2111,
        in1(1) => S2107,
        out1 => S2112
    );
nand_n_2685: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2108,
        in1(1) => S265,
        out1 => S2113
    );
nand_n_2686: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2113,
        in1(1) => S2112,
        out1 => S2114
    );
nand_n_2687: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2114,
        in1(1) => S2105,
        out1 => S2115
    );
nor_n_2688: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2083,
        in1(1) => S1995,
        out1 => S2116
    );
nand_n_2689: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2084,
        in1(1) => S1996,
        out1 => S2117
    );
nor_n_2690: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2022,
        in1(1) => S2001,
        out1 => S2118
    );
nand_n_2691: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2021,
        in1(1) => S2002,
        out1 => S2119
    );
nor_n_2692: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2118,
        in1(1) => S2023,
        out1 => S2120
    );
nand_n_2693: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2119,
        in1(1) => S2024,
        out1 => S2121
    );
nor_n_2694: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2120,
        in1(1) => S2084,
        out1 => S2122
    );
nand_n_2695: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2121,
        in1(1) => S2083,
        out1 => S2123
    );
nor_n_2696: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2122,
        in1(1) => S2116,
        out1 => S2124
    );
nand_n_2697: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2123,
        in1(1) => S2117,
        out1 => S2125
    );
nor_n_2698: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2124,
        in1(1) => S248,
        out1 => S2126
    );
nor_n_2699: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2104,
        in1(1) => S256,
        out1 => S2127
    );
nor_n_2700: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2127,
        in1(1) => S2126,
        out1 => S2128
    );
nand_n_2701: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2128,
        in1(1) => S2115,
        out1 => S2129
    );
nor_n_2702: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2125,
        in1(1) => S249,
        out1 => S2130
    );
nor_n_2703: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2083,
        in1(1) => S1981,
        out1 => S2131
    );
nand_n_2704: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2084,
        in1(1) => S1982,
        out1 => S2132
    );
nor_n_2705: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2026,
        in1(1) => S1987,
        out1 => S2133
    );
nand_n_2706: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2025,
        in1(1) => S1988,
        out1 => S2134
    );
nor_n_2707: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2133,
        in1(1) => S2027,
        out1 => S2135
    );
nand_n_2708: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2134,
        in1(1) => S2028,
        out1 => S2136
    );
nor_n_2709: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2135,
        in1(1) => S2084,
        out1 => S2137
    );
nand_n_2710: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2136,
        in1(1) => S2083,
        out1 => S2138
    );
nor_n_2711: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2137,
        in1(1) => S2131,
        out1 => S2139
    );
nand_n_2712: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2138,
        in1(1) => S2132,
        out1 => S2140
    );
nor_n_2713: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2140,
        in1(1) => S241,
        out1 => S2141
    );
nor_n_2714: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2141,
        in1(1) => S2130,
        out1 => S2142
    );
nand_n_2715: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2142,
        in1(1) => S2129,
        out1 => S2143
    );
nor_n_2716: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2098,
        in1(1) => S208,
        out1 => S2144
    );
nor_n_2717: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2139,
        in1(1) => S240,
        out1 => S2145
    );
nor_n_2718: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2145,
        in1(1) => S2144,
        out1 => S2146
    );
nand_n_2719: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2146,
        in1(1) => S2143,
        out1 => S2147
    );
nand_n_2720: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2147,
        in1(1) => S2099,
        out1 => S2148
    );
nand_n_2721: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2148,
        in1(1) => S2090,
        out1 => S2149
    );
nor_n_2722: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1953,
        in1(1) => S1952,
        out1 => S2150
    );
nor_n_2723: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2150,
        in1(1) => S2038,
        out1 => S2151
    );
notg_2724: ENTITY WORK.notg
    PORT MAP (
        in1 => S2151,
        out1 => S2152
    );
nand_n_2725: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2150,
        in1(1) => S2038,
        out1 => S2153
    );
notg_2726: ENTITY WORK.notg
    PORT MAP (
        in1 => S2153,
        out1 => S2154
    );
nor_n_2727: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2154,
        in1(1) => S2151,
        out1 => S2155
    );
nand_n_2728: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2153,
        in1(1) => S2152,
        out1 => S2156
    );
nor_n_2729: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2155,
        in1(1) => S2084,
        out1 => S2157
    );
nand_n_2730: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2156,
        in1(1) => S2083,
        out1 => S2158
    );
nor_n_2731: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2083,
        in1(1) => S1950,
        out1 => S2159
    );
nand_n_2732: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2084,
        in1(1) => S1951,
        out1 => S2160
    );
nor_n_2733: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2159,
        in1(1) => S2157,
        out1 => S2161
    );
nand_n_2734: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2160,
        in1(1) => S2158,
        out1 => S2162
    );
nor_n_2735: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2162,
        in1(1) => S229,
        out1 => S2163
    );
nor_n_2736: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2089,
        in1(1) => S203,
        out1 => S2164
    );
nor_n_2737: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2164,
        in1(1) => S2163,
        out1 => S2165
    );
nand_n_2738: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2165,
        in1(1) => S2149,
        out1 => S2166
    );
nor_n_2739: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2083,
        in1(1) => S1907,
        out1 => S2167
    );
nand_n_2740: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2084,
        in1(1) => S1906,
        out1 => S2168
    );
nand_n_2741: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1909,
        in1(1) => S1908,
        out1 => S2169
    );
nand_n_2742: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2169,
        in1(1) => S2053,
        out1 => S2170
    );
notg_2743: ENTITY WORK.notg
    PORT MAP (
        in1 => S2170,
        out1 => S2171
    );
nor_n_2744: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2169,
        in1(1) => S2053,
        out1 => S2172
    );
notg_2745: ENTITY WORK.notg
    PORT MAP (
        in1 => S2172,
        out1 => S2173
    );
nor_n_2746: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2172,
        in1(1) => S2171,
        out1 => S2174
    );
nand_n_2747: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2173,
        in1(1) => S2170,
        out1 => S2175
    );
nor_n_2748: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2175,
        in1(1) => S2084,
        out1 => S2176
    );
nand_n_2749: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2174,
        in1(1) => S2083,
        out1 => S2177
    );
nor_n_2750: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2176,
        in1(1) => S2167,
        out1 => S2178
    );
nand_n_2751: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2177,
        in1(1) => S2168,
        out1 => S2179
    );
nor_n_2752: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2178,
        in1(1) => new_datapath_multdivunit_1697_B_11,
        out1 => S2180
    );
nor_n_2753: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2179,
        in1(1) => S3445,
        out1 => S2181
    );
nor_n_2754: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2181,
        in1(1) => S2180,
        out1 => S2182
    );
nand_n_2755: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2049,
        in1(1) => S1919,
        out1 => S2183
    );
nand_n_2756: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2183,
        in1(1) => S2052,
        out1 => S2184
    );
nand_n_2757: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2184,
        in1(1) => S2083,
        out1 => S2185
    );
nand_n_2758: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2084,
        in1(1) => S1914,
        out1 => S2186
    );
nand_n_2759: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2186,
        in1(1) => S2185,
        out1 => S2187
    );
nor_n_2760: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2187,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S2188
    );
nand_n_2761: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2187,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S2189
    );
notg_2762: ENTITY WORK.notg
    PORT MAP (
        in1 => S2189,
        out1 => S2190
    );
nor_n_2763: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2190,
        in1(1) => S2188,
        out1 => S2191
    );
nand_n_2764: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2191,
        in1(1) => S2182,
        out1 => S2192
    );
nor_n_2765: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2161,
        in1(1) => S228,
        out1 => S2193
    );
nor_n_2766: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2042,
        in1(1) => S1942,
        out1 => S2194
    );
nor_n_2767: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2194,
        in1(1) => S2043,
        out1 => S2195
    );
nor_n_2768: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2195,
        in1(1) => S2084,
        out1 => S2196
    );
nor_n_2769: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2083,
        in1(1) => S1937,
        out1 => S2197
    );
nor_n_2770: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2197,
        in1(1) => S2196,
        out1 => S2198
    );
nor_n_2771: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2198,
        in1(1) => S3478,
        out1 => S2199
    );
nor_n_2772: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2199,
        in1(1) => S2193,
        out1 => S2200
    );
nand_n_2773: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1932,
        in1(1) => S1931,
        out1 => S2201
    );
nand_n_2774: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2201,
        in1(1) => S2045,
        out1 => S2202
    );
notg_2775: ENTITY WORK.notg
    PORT MAP (
        in1 => S2202,
        out1 => S2203
    );
nor_n_2776: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2201,
        in1(1) => S2045,
        out1 => S2204
    );
nor_n_2777: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2204,
        in1(1) => S2203,
        out1 => S2205
    );
nor_n_2778: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2205,
        in1(1) => S2084,
        out1 => S2206
    );
nor_n_2779: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2083,
        in1(1) => S1929,
        out1 => S2207
    );
nor_n_2780: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2207,
        in1(1) => S2206,
        out1 => S2208
    );
notg_2781: ENTITY WORK.notg
    PORT MAP (
        in1 => S2208,
        out1 => S2209
    );
nor_n_2782: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2208,
        in1(1) => S3467,
        out1 => S2210
    );
nand_n_2783: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2209,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S2211
    );
nand_n_2784: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2208,
        in1(1) => S3467,
        out1 => S2212
    );
nand_n_2785: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2198,
        in1(1) => S3478,
        out1 => S2213
    );
nand_n_2786: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2213,
        in1(1) => S2212,
        out1 => S2214
    );
nor_n_2787: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2214,
        in1(1) => S2210,
        out1 => S2215
    );
nand_n_2788: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2215,
        in1(1) => S2200,
        out1 => S2216
    );
nor_n_2789: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2216,
        in1(1) => S2192,
        out1 => S2217
    );
nand_n_2790: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2217,
        in1(1) => S2166,
        out1 => S2218
    );
nand_n_2791: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2214,
        in1(1) => S2211,
        out1 => S2219
    );
nor_n_2792: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2219,
        in1(1) => S2192,
        out1 => S2220
    );
nor_n_2793: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2188,
        in1(1) => S2180,
        out1 => S2221
    );
nor_n_2794: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2221,
        in1(1) => S2181,
        out1 => S2222
    );
nor_n_2795: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2222,
        in1(1) => S2220,
        out1 => S2223
    );
nand_n_2796: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2223,
        in1(1) => S2218,
        out1 => S2224
    );
nand_n_2797: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2065,
        in1(1) => S1867,
        out1 => S2225
    );
nand_n_2798: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2225,
        in1(1) => S2068,
        out1 => S2226
    );
nand_n_2799: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2226,
        in1(1) => S2083,
        out1 => S2227
    );
nand_n_2800: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2084,
        in1(1) => S1862,
        out1 => S2228
    );
nand_n_2801: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2228,
        in1(1) => S2227,
        out1 => S2229
    );
nand_n_2802: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2069,
        in1(1) => S3412,
        out1 => S2230
    );
notg_2803: ENTITY WORK.notg
    PORT MAP (
        in1 => S2230,
        out1 => S2231
    );
nand_n_2804: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1848,
        in1(1) => new_datapath_multdivunit_1697_B_15,
        out1 => S2232
    );
nand_n_2805: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2229,
        in1(1) => new_datapath_multdivunit_1697_B_14,
        out1 => S2233
    );
notg_2806: ENTITY WORK.notg
    PORT MAP (
        in1 => S2233,
        out1 => S2234
    );
nor_n_2807: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2229,
        in1(1) => new_datapath_multdivunit_1697_B_14,
        out1 => S2235
    );
nor_n_2808: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2069,
        in1(1) => S3412,
        out1 => S2236
    );
nor_n_2809: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2236,
        in1(1) => S2231,
        out1 => S2237
    );
nand_n_2810: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2237,
        in1(1) => S2080,
        out1 => S2238
    );
nor_n_2811: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2235,
        in1(1) => S2234,
        out1 => S2239
    );
nand_n_2812: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2238,
        in1(1) => S2232,
        out1 => S2240
    );
notg_2813: ENTITY WORK.notg
    PORT MAP (
        in1 => S2240,
        out1 => S2241
    );
nand_n_2814: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2241,
        in1(1) => S2239,
        out1 => S2242
    );
nand_n_2815: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1881,
        in1(1) => S1880,
        out1 => S2243
    );
nand_n_2816: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2243,
        in1(1) => S2061,
        out1 => S2244
    );
notg_2817: ENTITY WORK.notg
    PORT MAP (
        in1 => S2244,
        out1 => S2245
    );
nor_n_2818: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2243,
        in1(1) => S2061,
        out1 => S2246
    );
notg_2819: ENTITY WORK.notg
    PORT MAP (
        in1 => S2246,
        out1 => S2247
    );
nor_n_2820: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2246,
        in1(1) => S2245,
        out1 => S2248
    );
nand_n_2821: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2247,
        in1(1) => S2244,
        out1 => S2249
    );
nor_n_2822: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2248,
        in1(1) => S2084,
        out1 => S2250
    );
nand_n_2823: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2249,
        in1(1) => S2083,
        out1 => S2251
    );
nor_n_2824: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2083,
        in1(1) => S1878,
        out1 => S2252
    );
nand_n_2825: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2084,
        in1(1) => S1879,
        out1 => S2253
    );
nor_n_2826: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2252,
        in1(1) => S2250,
        out1 => S2254
    );
nand_n_2827: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2253,
        in1(1) => S2251,
        out1 => S2255
    );
nor_n_2828: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2255,
        in1(1) => new_datapath_multdivunit_1697_B_13,
        out1 => S2256
    );
nand_n_2829: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2254,
        in1(1) => S3423,
        out1 => S2257
    );
nor_n_2830: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2058,
        in1(1) => S1895,
        out1 => S2258
    );
nor_n_2831: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2258,
        in1(1) => S2059,
        out1 => S2259
    );
nor_n_2832: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2259,
        in1(1) => S2084,
        out1 => S2260
    );
nor_n_2833: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2083,
        in1(1) => S1889,
        out1 => S2261
    );
nor_n_2834: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2261,
        in1(1) => S2260,
        out1 => S2262
    );
notg_2835: ENTITY WORK.notg
    PORT MAP (
        in1 => S2262,
        out1 => S2263
    );
nor_n_2836: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2263,
        in1(1) => new_datapath_multdivunit_1697_B_12,
        out1 => S2264
    );
nand_n_2837: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2262,
        in1(1) => S3434,
        out1 => S2265
    );
nor_n_2838: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2264,
        in1(1) => S2256,
        out1 => S2266
    );
nand_n_2839: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2265,
        in1(1) => S2257,
        out1 => S2267
    );
nor_n_2840: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2254,
        in1(1) => S3423,
        out1 => S2268
    );
nand_n_2841: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2255,
        in1(1) => new_datapath_multdivunit_1697_B_13,
        out1 => S2269
    );
nor_n_2842: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2262,
        in1(1) => S3434,
        out1 => S2270
    );
nor_n_2843: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2270,
        in1(1) => S2268,
        out1 => S2271
    );
nand_n_2844: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2271,
        in1(1) => S2266,
        out1 => S2272
    );
nor_n_2845: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2272,
        in1(1) => S2242,
        out1 => S2273
    );
nand_n_2846: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2273,
        in1(1) => S2224,
        out1 => S2274
    );
nand_n_2847: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2269,
        in1(1) => S2267,
        out1 => S2275
    );
nor_n_2848: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2275,
        in1(1) => S2242,
        out1 => S2276
    );
nand_n_2849: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2235,
        in1(1) => S2232,
        out1 => S2277
    );
nand_n_2850: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2277,
        in1(1) => S2238,
        out1 => S2278
    );
nor_n_2851: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2278,
        in1(1) => S2276,
        out1 => S2279
    );
nand_n_2852: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2279,
        in1(1) => S2274,
        out1 => S2280
    );
nand_n_2853: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2280,
        in1(1) => S5537,
        out1 => S2281
    );
nand_n_2854: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5611,
        in1(1) => new_datapath_multdivunit_outmdu1_0,
        out1 => S2282
    );
nor_n_2855: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => S5590,
        out1 => S2283
    );
nand_n_2856: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2283,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S2284
    );
nand_n_2857: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2284,
        in1(1) => S2282,
        out1 => S2285
    );
notg_2858: ENTITY WORK.notg
    PORT MAP (
        in1 => S2285,
        out1 => S2286
    );
nand_n_2859: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2286,
        in1(1) => S2281,
        out1 => S20
    );
nor_n_2860: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2084,
        in1(1) => S5547,
        out1 => S2287
    );
nand_n_2861: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5611,
        in1(1) => new_datapath_multdivunit_outmdu1_1,
        out1 => S2288
    );
nor_n_2862: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => S5966,
        out1 => S2289
    );
nor_n_2863: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S264,
        in1(1) => S5975,
        out1 => S2290
    );
nand_n_2864: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S265,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S2291
    );
nand_n_2865: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2290,
        in1(1) => S2289,
        out1 => S2292
    );
nor_n_2866: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2290,
        in1(1) => S2289,
        out1 => S2293
    );
nand_n_2867: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2292,
        in1(1) => S5579,
        out1 => S2294
    );
nor_n_2868: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2294,
        in1(1) => S2293,
        out1 => S2295
    );
nor_n_2869: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2295,
        in1(1) => S2287,
        out1 => S2296
    );
nand_n_2870: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2296,
        in1(1) => S2288,
        out1 => S21
    );
nor_n_2871: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1857,
        in1(1) => S5547,
        out1 => S2297
    );
nor_n_2872: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S256,
        in1(1) => S5975,
        out1 => S2298
    );
nand_n_2873: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S2299
    );
nand_n_2874: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S2300
    );
nand_n_2875: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2300,
        in1(1) => S2291,
        out1 => S2301
    );
nor_n_2876: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S264,
        in1(1) => S5957,
        out1 => S2302
    );
nand_n_2877: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S265,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S2303
    );
nand_n_2878: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2302,
        in1(1) => S2289,
        out1 => S2304
    );
nand_n_2879: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2304,
        in1(1) => S2301,
        out1 => S2305
    );
notg_2880: ENTITY WORK.notg
    PORT MAP (
        in1 => S2305,
        out1 => S2306
    );
nand_n_2881: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2306,
        in1(1) => S2298,
        out1 => S2307
    );
nand_n_2882: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2305,
        in1(1) => S2299,
        out1 => S2308
    );
nand_n_2883: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2308,
        in1(1) => S2307,
        out1 => S2309
    );
nand_n_2884: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2309,
        in1(1) => S2292,
        out1 => S2310
    );
nor_n_2885: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2309,
        in1(1) => S2292,
        out1 => S2311
    );
nor_n_2886: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2311,
        in1(1) => S5590,
        out1 => S2312
    );
nand_n_2887: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2312,
        in1(1) => S2310,
        out1 => S2313
    );
nand_n_2888: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5611,
        in1(1) => new_datapath_multdivunit_outmdu1_2,
        out1 => S2314
    );
notg_2889: ENTITY WORK.notg
    PORT MAP (
        in1 => S2314,
        out1 => S2315
    );
nor_n_2890: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2315,
        in1(1) => S2297,
        out1 => S2316
    );
nand_n_2891: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2316,
        in1(1) => S2313,
        out1 => S22
    );
nor_n_2892: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1635,
        in1(1) => S5547,
        out1 => S2317
    );
nand_n_2893: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5611,
        in1(1) => new_datapath_multdivunit_outmdu1_3,
        out1 => S2318
    );
nor_n_2894: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S248,
        in1(1) => S5975,
        out1 => S2319
    );
nand_n_2895: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S249,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S2320
    );
nand_n_2896: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2307,
        in1(1) => S2304,
        out1 => S2321
    );
notg_2897: ENTITY WORK.notg
    PORT MAP (
        in1 => S2321,
        out1 => S2322
    );
nor_n_2898: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S256,
        in1(1) => S5966,
        out1 => S2323
    );
nand_n_2899: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S2324
    );
nor_n_2900: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => S5947,
        out1 => S2325
    );
nand_n_2901: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S2326
    );
nor_n_2902: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2325,
        in1(1) => S2302,
        out1 => S2327
    );
nand_n_2903: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2326,
        in1(1) => S2303,
        out1 => S2328
    );
nor_n_2904: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S264,
        in1(1) => S5947,
        out1 => S2329
    );
nand_n_2905: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S265,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S2330
    );
nor_n_2906: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2326,
        in1(1) => S2303,
        out1 => S2331
    );
nand_n_2907: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2325,
        in1(1) => S2302,
        out1 => S2332
    );
nor_n_2908: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2331,
        in1(1) => S2327,
        out1 => S2333
    );
nand_n_2909: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2332,
        in1(1) => S2328,
        out1 => S2334
    );
nor_n_2910: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2334,
        in1(1) => S2324,
        out1 => S2335
    );
nand_n_2911: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2333,
        in1(1) => S2323,
        out1 => S2336
    );
nor_n_2912: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2333,
        in1(1) => S2323,
        out1 => S2337
    );
nand_n_2913: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2334,
        in1(1) => S2324,
        out1 => S2338
    );
nor_n_2914: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2337,
        in1(1) => S2335,
        out1 => S2339
    );
nand_n_2915: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2338,
        in1(1) => S2336,
        out1 => S2340
    );
nor_n_2916: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2340,
        in1(1) => S2322,
        out1 => S2341
    );
nor_n_2917: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2339,
        in1(1) => S2321,
        out1 => S2342
    );
nor_n_2918: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2342,
        in1(1) => S2341,
        out1 => S2343
    );
notg_2919: ENTITY WORK.notg
    PORT MAP (
        in1 => S2343,
        out1 => S2344
    );
nor_n_2920: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2344,
        in1(1) => S2320,
        out1 => S2345
    );
nor_n_2921: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2343,
        in1(1) => S2319,
        out1 => S2346
    );
nor_n_2922: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2346,
        in1(1) => S2345,
        out1 => S2347
    );
nand_n_2923: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2347,
        in1(1) => S2311,
        out1 => S2348
    );
nor_n_2924: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2347,
        in1(1) => S2311,
        out1 => S2349
    );
nand_n_2925: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2348,
        in1(1) => S5579,
        out1 => S2350
    );
nor_n_2926: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2350,
        in1(1) => S2349,
        out1 => S2351
    );
nor_n_2927: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2351,
        in1(1) => S2317,
        out1 => S2352
    );
nand_n_2928: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2352,
        in1(1) => S2318,
        out1 => S23
    );
nor_n_2929: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S1452,
        in1(1) => S5547,
        out1 => S2353
    );
nand_n_2930: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5611,
        in1(1) => new_datapath_multdivunit_outmdu1_4,
        out1 => S2354
    );
nor_n_2931: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2345,
        in1(1) => S2341,
        out1 => S2355
    );
notg_2932: ENTITY WORK.notg
    PORT MAP (
        in1 => S2355,
        out1 => S2356
    );
nand_n_2933: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S241,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S2357
    );
nand_n_2934: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S249,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S2358
    );
nand_n_2935: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2358,
        in1(1) => S2357,
        out1 => S2359
    );
nor_n_2936: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S240,
        in1(1) => S5966,
        out1 => S2360
    );
nand_n_2937: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S241,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S2361
    );
nor_n_2938: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2361,
        in1(1) => S2320,
        out1 => S2362
    );
nand_n_2939: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2360,
        in1(1) => S2319,
        out1 => S2363
    );
nand_n_2940: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2363,
        in1(1) => S2359,
        out1 => S2364
    );
notg_2941: ENTITY WORK.notg
    PORT MAP (
        in1 => S2364,
        out1 => S2365
    );
nor_n_2942: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2335,
        in1(1) => S2331,
        out1 => S2366
    );
nand_n_2943: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2336,
        in1(1) => S2332,
        out1 => S2367
    );
nor_n_2944: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S256,
        in1(1) => S5957,
        out1 => S2368
    );
nand_n_2945: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S2369
    );
nor_n_2946: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2329,
        in1(1) => S1204,
        out1 => S2370
    );
nand_n_2947: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2330,
        in1(1) => S1205,
        out1 => S2371
    );
nor_n_2948: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S264,
        in1(1) => S5936,
        out1 => S2372
    );
nand_n_2949: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S265,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S2373
    );
nor_n_2950: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2330,
        in1(1) => S1205,
        out1 => S2374
    );
nand_n_2951: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2329,
        in1(1) => S1204,
        out1 => S2375
    );
nor_n_2952: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2374,
        in1(1) => S2370,
        out1 => S2376
    );
nand_n_2953: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2375,
        in1(1) => S2371,
        out1 => S2377
    );
nor_n_2954: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2377,
        in1(1) => S2369,
        out1 => S2378
    );
nand_n_2955: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2376,
        in1(1) => S2368,
        out1 => S2379
    );
nor_n_2956: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2376,
        in1(1) => S2368,
        out1 => S2380
    );
nand_n_2957: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2377,
        in1(1) => S2369,
        out1 => S2381
    );
nor_n_2958: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2380,
        in1(1) => S2378,
        out1 => S2382
    );
nand_n_2959: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2381,
        in1(1) => S2379,
        out1 => S2383
    );
nor_n_2960: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2383,
        in1(1) => S2366,
        out1 => S2384
    );
nand_n_2961: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2382,
        in1(1) => S2367,
        out1 => S2385
    );
nand_n_2962: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2383,
        in1(1) => S2366,
        out1 => S2386
    );
nand_n_2963: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2386,
        in1(1) => S2385,
        out1 => S2387
    );
notg_2964: ENTITY WORK.notg
    PORT MAP (
        in1 => S2387,
        out1 => S2388
    );
nand_n_2965: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2388,
        in1(1) => S2365,
        out1 => S2389
    );
notg_2966: ENTITY WORK.notg
    PORT MAP (
        in1 => S2389,
        out1 => S2390
    );
nand_n_2967: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2387,
        in1(1) => S2364,
        out1 => S2391
    );
nand_n_2968: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2391,
        in1(1) => S2389,
        out1 => S2392
    );
notg_2969: ENTITY WORK.notg
    PORT MAP (
        in1 => S2392,
        out1 => S2393
    );
nand_n_2970: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2392,
        in1(1) => S2355,
        out1 => S2394
    );
nand_n_2971: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2393,
        in1(1) => S2356,
        out1 => S2395
    );
notg_2972: ENTITY WORK.notg
    PORT MAP (
        in1 => S2395,
        out1 => S2396
    );
nand_n_2973: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2395,
        in1(1) => S2394,
        out1 => S2397
    );
nor_n_2974: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2397,
        in1(1) => S2348,
        out1 => S2398
    );
notg_2975: ENTITY WORK.notg
    PORT MAP (
        in1 => S2398,
        out1 => S2399
    );
nand_n_2976: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2397,
        in1(1) => S2348,
        out1 => S2400
    );
nand_n_2977: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2400,
        in1(1) => S5579,
        out1 => S2401
    );
nor_n_2978: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2401,
        in1(1) => S2398,
        out1 => S2402
    );
nor_n_2979: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2402,
        in1(1) => S2353,
        out1 => S2403
    );
nand_n_2980: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2403,
        in1(1) => S2354,
        out1 => S24
    );
nand_n_2981: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1267,
        in1(1) => S5537,
        out1 => S2404
    );
nor_n_2982: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2390,
        in1(1) => S2384,
        out1 => S2405
    );
nand_n_2983: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2389,
        in1(1) => S2385,
        out1 => S2406
    );
nor_n_2984: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S208,
        in1(1) => S5975,
        out1 => S2407
    );
nand_n_2985: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S209,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S2408
    );
nor_n_2986: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S248,
        in1(1) => S5957,
        out1 => S2409
    );
nand_n_2987: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S249,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S2410
    );
nor_n_2988: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2409,
        in1(1) => S2360,
        out1 => S2411
    );
nand_n_2989: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2410,
        in1(1) => S2361,
        out1 => S2412
    );
nor_n_2990: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S240,
        in1(1) => S5957,
        out1 => S2413
    );
nand_n_2991: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S241,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S2414
    );
nor_n_2992: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2410,
        in1(1) => S2361,
        out1 => S2415
    );
nand_n_2993: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2409,
        in1(1) => S2360,
        out1 => S2416
    );
nor_n_2994: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2415,
        in1(1) => S2411,
        out1 => S2417
    );
nand_n_2995: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2416,
        in1(1) => S2412,
        out1 => S2418
    );
nor_n_2996: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2418,
        in1(1) => S2408,
        out1 => S2419
    );
nand_n_2997: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2417,
        in1(1) => S2407,
        out1 => S2420
    );
nor_n_2998: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2417,
        in1(1) => S2407,
        out1 => S2421
    );
nand_n_2999: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2418,
        in1(1) => S2408,
        out1 => S2422
    );
nor_n_3000: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2421,
        in1(1) => S2419,
        out1 => S2423
    );
nand_n_3001: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2422,
        in1(1) => S2420,
        out1 => S2424
    );
nor_n_3002: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2378,
        in1(1) => S2374,
        out1 => S2425
    );
nand_n_3003: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2379,
        in1(1) => S2375,
        out1 => S2426
    );
nor_n_3004: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S256,
        in1(1) => S5947,
        out1 => S2427
    );
nand_n_3005: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S2428
    );
nor_n_3006: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2372,
        in1(1) => S1208,
        out1 => S2429
    );
nand_n_3007: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2373,
        in1(1) => S1209,
        out1 => S2430
    );
nor_n_3008: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S264,
        in1(1) => S5926,
        out1 => S2431
    );
nand_n_3009: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S265,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S2432
    );
nor_n_3010: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2373,
        in1(1) => S1209,
        out1 => S2433
    );
nand_n_3011: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2372,
        in1(1) => S1208,
        out1 => S2434
    );
nor_n_3012: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2433,
        in1(1) => S2429,
        out1 => S2435
    );
nand_n_3013: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2434,
        in1(1) => S2430,
        out1 => S2436
    );
nor_n_3014: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2436,
        in1(1) => S2428,
        out1 => S2437
    );
nand_n_3015: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2435,
        in1(1) => S2427,
        out1 => S2438
    );
nor_n_3016: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2435,
        in1(1) => S2427,
        out1 => S2439
    );
nand_n_3017: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2436,
        in1(1) => S2428,
        out1 => S2440
    );
nor_n_3018: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2439,
        in1(1) => S2437,
        out1 => S2441
    );
nand_n_3019: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2440,
        in1(1) => S2438,
        out1 => S2442
    );
nor_n_3020: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2442,
        in1(1) => S2425,
        out1 => S2443
    );
nand_n_3021: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2441,
        in1(1) => S2426,
        out1 => S2444
    );
nor_n_3022: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2441,
        in1(1) => S2426,
        out1 => S2445
    );
nand_n_3023: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2442,
        in1(1) => S2425,
        out1 => S2446
    );
nor_n_3024: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2445,
        in1(1) => S2443,
        out1 => S2447
    );
nand_n_3025: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2446,
        in1(1) => S2444,
        out1 => S2448
    );
nor_n_3026: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2448,
        in1(1) => S2424,
        out1 => S2449
    );
nand_n_3027: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2447,
        in1(1) => S2423,
        out1 => S2450
    );
nor_n_3028: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2447,
        in1(1) => S2423,
        out1 => S2451
    );
nand_n_3029: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2448,
        in1(1) => S2424,
        out1 => S2452
    );
nor_n_3030: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2451,
        in1(1) => S2449,
        out1 => S2453
    );
nand_n_3031: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2452,
        in1(1) => S2450,
        out1 => S2454
    );
nand_n_3032: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2453,
        in1(1) => S2406,
        out1 => S2455
    );
nand_n_3033: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2454,
        in1(1) => S2405,
        out1 => S2456
    );
nand_n_3034: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2456,
        in1(1) => S2455,
        out1 => S2457
    );
notg_3035: ENTITY WORK.notg
    PORT MAP (
        in1 => S2457,
        out1 => S2458
    );
nand_n_3036: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2458,
        in1(1) => S2362,
        out1 => S2459
    );
nand_n_3037: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2457,
        in1(1) => S2363,
        out1 => S2460
    );
nand_n_3038: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2460,
        in1(1) => S2459,
        out1 => S2461
    );
notg_3039: ENTITY WORK.notg
    PORT MAP (
        in1 => S2461,
        out1 => S2462
    );
nand_n_3040: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2462,
        in1(1) => S2396,
        out1 => S2463
    );
nand_n_3041: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2461,
        in1(1) => S2395,
        out1 => S2464
    );
nand_n_3042: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2464,
        in1(1) => S2463,
        out1 => S2465
    );
nor_n_3043: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2465,
        in1(1) => S2399,
        out1 => S2466
    );
notg_3044: ENTITY WORK.notg
    PORT MAP (
        in1 => S2466,
        out1 => S2467
    );
nand_n_3045: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2465,
        in1(1) => S2399,
        out1 => S2468
    );
nand_n_3046: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2468,
        in1(1) => S5579,
        out1 => S2469
    );
nor_n_3047: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2469,
        in1(1) => S2466,
        out1 => S2470
    );
nand_n_3048: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5611,
        in1(1) => new_datapath_multdivunit_outmdu1_5,
        out1 => S2471
    );
notg_3049: ENTITY WORK.notg
    PORT MAP (
        in1 => S2471,
        out1 => S2472
    );
nor_n_3050: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2472,
        in1(1) => S2470,
        out1 => S2473
    );
nand_n_3051: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2473,
        in1(1) => S2404,
        out1 => S25
    );
nand_n_3052: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S1084,
        in1(1) => S5537,
        out1 => S2474
    );
nor_n_3053: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5600,
        in1(1) => S2789,
        out1 => S2475
    );
nand_n_3054: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2459,
        in1(1) => S2455,
        out1 => S2476
    );
notg_3055: ENTITY WORK.notg
    PORT MAP (
        in1 => S2476,
        out1 => S2477
    );
nor_n_3056: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S202,
        in1(1) => S5975,
        out1 => S2478
    );
nand_n_3057: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S203,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S2479
    );
nor_n_3058: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2419,
        in1(1) => S2415,
        out1 => S2480
    );
nand_n_3059: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2420,
        in1(1) => S2416,
        out1 => S2481
    );
nor_n_3060: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2480,
        in1(1) => S2479,
        out1 => S2482
    );
nand_n_3061: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2481,
        in1(1) => S2478,
        out1 => S2483
    );
nor_n_3062: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2481,
        in1(1) => S2478,
        out1 => S2484
    );
nand_n_3063: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2480,
        in1(1) => S2479,
        out1 => S2485
    );
nor_n_3064: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2484,
        in1(1) => S2482,
        out1 => S2486
    );
nand_n_3065: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2485,
        in1(1) => S2483,
        out1 => S2487
    );
nor_n_3066: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2449,
        in1(1) => S2443,
        out1 => S2488
    );
nand_n_3067: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2450,
        in1(1) => S2444,
        out1 => S2489
    );
nor_n_3068: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S208,
        in1(1) => S5966,
        out1 => S2490
    );
nand_n_3069: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S209,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S2491
    );
nor_n_3070: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S248,
        in1(1) => S5947,
        out1 => S2492
    );
nand_n_3071: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S249,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S2493
    );
nor_n_3072: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2492,
        in1(1) => S2413,
        out1 => S2494
    );
nand_n_3073: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2493,
        in1(1) => S2414,
        out1 => S2495
    );
nor_n_3074: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S240,
        in1(1) => S5947,
        out1 => S2496
    );
nand_n_3075: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S241,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S2497
    );
nor_n_3076: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2493,
        in1(1) => S2414,
        out1 => S2498
    );
nand_n_3077: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2492,
        in1(1) => S2413,
        out1 => S2499
    );
nor_n_3078: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2498,
        in1(1) => S2494,
        out1 => S2500
    );
nand_n_3079: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2499,
        in1(1) => S2495,
        out1 => S2501
    );
nor_n_3080: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2501,
        in1(1) => S2491,
        out1 => S2502
    );
nand_n_3081: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2500,
        in1(1) => S2490,
        out1 => S2503
    );
nor_n_3082: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2500,
        in1(1) => S2490,
        out1 => S2504
    );
nand_n_3083: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2501,
        in1(1) => S2491,
        out1 => S2505
    );
nor_n_3084: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2504,
        in1(1) => S2502,
        out1 => S2506
    );
nand_n_3085: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2505,
        in1(1) => S2503,
        out1 => S2507
    );
nor_n_3086: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2437,
        in1(1) => S2433,
        out1 => S2508
    );
nand_n_3087: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2438,
        in1(1) => S2434,
        out1 => S2509
    );
nor_n_3088: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S256,
        in1(1) => S5936,
        out1 => S2510
    );
nand_n_3089: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S2511
    );
nor_n_3090: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2431,
        in1(1) => S882,
        out1 => S2512
    );
nand_n_3091: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2432,
        in1(1) => S883,
        out1 => S2513
    );
nor_n_3092: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S264,
        in1(1) => S5916,
        out1 => S2514
    );
nand_n_3093: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S265,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S2515
    );
nor_n_3094: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2432,
        in1(1) => S883,
        out1 => S2516
    );
nand_n_3095: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2431,
        in1(1) => S882,
        out1 => S2517
    );
nor_n_3096: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2516,
        in1(1) => S2512,
        out1 => S2518
    );
nand_n_3097: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2517,
        in1(1) => S2513,
        out1 => S2519
    );
nor_n_3098: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2519,
        in1(1) => S2511,
        out1 => S2520
    );
nand_n_3099: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2518,
        in1(1) => S2510,
        out1 => S2521
    );
nor_n_3100: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2518,
        in1(1) => S2510,
        out1 => S2522
    );
nand_n_3101: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2519,
        in1(1) => S2511,
        out1 => S2523
    );
nor_n_3102: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2522,
        in1(1) => S2520,
        out1 => S2524
    );
nand_n_3103: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2523,
        in1(1) => S2521,
        out1 => S2525
    );
nor_n_3104: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2525,
        in1(1) => S2508,
        out1 => S2526
    );
nand_n_3105: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2524,
        in1(1) => S2509,
        out1 => S2527
    );
nor_n_3106: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2524,
        in1(1) => S2509,
        out1 => S2528
    );
nand_n_3107: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2525,
        in1(1) => S2508,
        out1 => S2529
    );
nor_n_3108: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2528,
        in1(1) => S2526,
        out1 => S2530
    );
nand_n_3109: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2529,
        in1(1) => S2527,
        out1 => S2531
    );
nor_n_3110: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2531,
        in1(1) => S2507,
        out1 => S2532
    );
nand_n_3111: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2530,
        in1(1) => S2506,
        out1 => S2533
    );
nor_n_3112: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2530,
        in1(1) => S2506,
        out1 => S2534
    );
nand_n_3113: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2531,
        in1(1) => S2507,
        out1 => S2535
    );
nor_n_3114: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2534,
        in1(1) => S2532,
        out1 => S2536
    );
nand_n_3115: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2535,
        in1(1) => S2533,
        out1 => S2537
    );
nor_n_3116: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2537,
        in1(1) => S2488,
        out1 => S2538
    );
nand_n_3117: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2536,
        in1(1) => S2489,
        out1 => S2539
    );
nor_n_3118: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2536,
        in1(1) => S2489,
        out1 => S2540
    );
nand_n_3119: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2537,
        in1(1) => S2488,
        out1 => S2541
    );
nor_n_3120: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2540,
        in1(1) => S2538,
        out1 => S2542
    );
nand_n_3121: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2541,
        in1(1) => S2539,
        out1 => S2543
    );
nor_n_3122: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2543,
        in1(1) => S2487,
        out1 => S2544
    );
nand_n_3123: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2542,
        in1(1) => S2486,
        out1 => S2545
    );
nor_n_3124: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2542,
        in1(1) => S2486,
        out1 => S2546
    );
nand_n_3125: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2543,
        in1(1) => S2487,
        out1 => S2547
    );
nor_n_3126: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2546,
        in1(1) => S2544,
        out1 => S2548
    );
nand_n_3127: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2547,
        in1(1) => S2545,
        out1 => S2549
    );
nand_n_3128: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2549,
        in1(1) => S2477,
        out1 => S2550
    );
nand_n_3129: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2548,
        in1(1) => S2476,
        out1 => S2551
    );
notg_3130: ENTITY WORK.notg
    PORT MAP (
        in1 => S2551,
        out1 => S2552
    );
nand_n_3131: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2551,
        in1(1) => S2550,
        out1 => S2553
    );
nor_n_3132: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2553,
        in1(1) => S2463,
        out1 => S2554
    );
nand_n_3133: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2553,
        in1(1) => S2463,
        out1 => S2555
    );
notg_3134: ENTITY WORK.notg
    PORT MAP (
        in1 => S2555,
        out1 => S2556
    );
nor_n_3135: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2556,
        in1(1) => S2554,
        out1 => S2557
    );
notg_3136: ENTITY WORK.notg
    PORT MAP (
        in1 => S2557,
        out1 => S2558
    );
nor_n_3137: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2558,
        in1(1) => S2467,
        out1 => S2559
    );
nand_n_3138: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2558,
        in1(1) => S2467,
        out1 => S2560
    );
nand_n_3139: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2560,
        in1(1) => S5579,
        out1 => S2561
    );
nor_n_3140: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2561,
        in1(1) => S2559,
        out1 => S2562
    );
nor_n_3141: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2562,
        in1(1) => S2475,
        out1 => S2563
    );
nand_n_3142: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2563,
        in1(1) => S2474,
        out1 => S26
    );
nor_n_3143: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S937,
        in1(1) => S5547,
        out1 => S2564
    );
nand_n_3144: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5611,
        in1(1) => new_datapath_multdivunit_outmdu1_7,
        out1 => S2565
    );
nor_n_3145: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2544,
        in1(1) => S2538,
        out1 => S2566
    );
nand_n_3146: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2545,
        in1(1) => S2539,
        out1 => S2567
    );
nor_n_3147: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S228,
        in1(1) => S5975,
        out1 => S2568
    );
nand_n_3148: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S229,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S2569
    );
nor_n_3149: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S202,
        in1(1) => S5966,
        out1 => S2570
    );
nand_n_3150: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S203,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S2571
    );
nor_n_3151: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2570,
        in1(1) => S2568,
        out1 => S2572
    );
nand_n_3152: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2571,
        in1(1) => S2569,
        out1 => S2573
    );
nor_n_3153: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S228,
        in1(1) => S5966,
        out1 => S2574
    );
nand_n_3154: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S229,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S2575
    );
nor_n_3155: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2575,
        in1(1) => S2479,
        out1 => S2576
    );
nand_n_3156: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2574,
        in1(1) => S2478,
        out1 => S2577
    );
nor_n_3157: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2576,
        in1(1) => S2572,
        out1 => S2578
    );
nand_n_3158: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2577,
        in1(1) => S2573,
        out1 => S2579
    );
nor_n_3159: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2502,
        in1(1) => S2498,
        out1 => S2580
    );
nand_n_3160: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2503,
        in1(1) => S2499,
        out1 => S2582
    );
nor_n_3161: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2582,
        in1(1) => S2578,
        out1 => S2583
    );
nand_n_3162: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2580,
        in1(1) => S2579,
        out1 => S2584
    );
nor_n_3163: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2580,
        in1(1) => S2579,
        out1 => S2585
    );
nand_n_3164: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2582,
        in1(1) => S2578,
        out1 => S2586
    );
nor_n_3165: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2585,
        in1(1) => S2583,
        out1 => S2587
    );
nand_n_3166: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2586,
        in1(1) => S2584,
        out1 => S2588
    );
nor_n_3167: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2532,
        in1(1) => S2526,
        out1 => S2589
    );
nand_n_3168: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2533,
        in1(1) => S2527,
        out1 => S2590
    );
nor_n_3169: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S208,
        in1(1) => S5957,
        out1 => S2591
    );
nand_n_3170: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S209,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S2593
    );
nor_n_3171: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S248,
        in1(1) => S5936,
        out1 => S2594
    );
nand_n_3172: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S249,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S2595
    );
nor_n_3173: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2594,
        in1(1) => S2496,
        out1 => S2596
    );
nand_n_3174: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2595,
        in1(1) => S2497,
        out1 => S2597
    );
nor_n_3175: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S240,
        in1(1) => S5936,
        out1 => S2598
    );
nand_n_3176: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S241,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S2599
    );
nor_n_3177: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2595,
        in1(1) => S2497,
        out1 => S2600
    );
nand_n_3178: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2594,
        in1(1) => S2496,
        out1 => S2601
    );
nor_n_3179: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2600,
        in1(1) => S2596,
        out1 => S2602
    );
nand_n_3180: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2601,
        in1(1) => S2597,
        out1 => S2604
    );
nor_n_3181: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2604,
        in1(1) => S2593,
        out1 => S2605
    );
nand_n_3182: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2602,
        in1(1) => S2591,
        out1 => S2606
    );
nor_n_3183: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2602,
        in1(1) => S2591,
        out1 => S2607
    );
nand_n_3184: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2604,
        in1(1) => S2593,
        out1 => S2608
    );
nor_n_3185: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2607,
        in1(1) => S2605,
        out1 => S2609
    );
nand_n_3186: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2608,
        in1(1) => S2606,
        out1 => S2610
    );
nor_n_3187: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2520,
        in1(1) => S2516,
        out1 => S2611
    );
nand_n_3188: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2521,
        in1(1) => S2517,
        out1 => S2612
    );
nor_n_3189: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S256,
        in1(1) => S5926,
        out1 => S2613
    );
nand_n_3190: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S2615
    );
nor_n_3191: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2514,
        in1(1) => S886,
        out1 => S2616
    );
nand_n_3192: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2515,
        in1(1) => S887,
        out1 => S2617
    );
nand_n_3193: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S265,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S2618
    );
nor_n_3194: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2515,
        in1(1) => S887,
        out1 => S2619
    );
nand_n_3195: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2514,
        in1(1) => S886,
        out1 => S2620
    );
nor_n_3196: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2619,
        in1(1) => S2616,
        out1 => S2621
    );
nand_n_3197: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2620,
        in1(1) => S2617,
        out1 => S2622
    );
nor_n_3198: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2622,
        in1(1) => S2615,
        out1 => S2623
    );
nand_n_3199: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2621,
        in1(1) => S2613,
        out1 => S2624
    );
nor_n_3200: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2621,
        in1(1) => S2613,
        out1 => S2626
    );
nand_n_3201: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2622,
        in1(1) => S2615,
        out1 => S2627
    );
nor_n_3202: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2626,
        in1(1) => S2623,
        out1 => S2628
    );
nand_n_3203: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2627,
        in1(1) => S2624,
        out1 => S2629
    );
nor_n_3204: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2629,
        in1(1) => S2611,
        out1 => S2630
    );
nand_n_3205: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2628,
        in1(1) => S2612,
        out1 => S2631
    );
nor_n_3206: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2628,
        in1(1) => S2612,
        out1 => S2632
    );
nand_n_3207: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2629,
        in1(1) => S2611,
        out1 => S2633
    );
nor_n_3208: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2632,
        in1(1) => S2630,
        out1 => S2634
    );
nand_n_3209: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2633,
        in1(1) => S2631,
        out1 => S2635
    );
nor_n_3210: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2635,
        in1(1) => S2610,
        out1 => S2637
    );
nand_n_3211: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2634,
        in1(1) => S2609,
        out1 => S2638
    );
nor_n_3212: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2634,
        in1(1) => S2609,
        out1 => S2639
    );
nand_n_3213: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2635,
        in1(1) => S2610,
        out1 => S2640
    );
nor_n_3214: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2639,
        in1(1) => S2637,
        out1 => S2641
    );
nand_n_3215: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2640,
        in1(1) => S2638,
        out1 => S2642
    );
nor_n_3216: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2642,
        in1(1) => S2589,
        out1 => S2643
    );
nand_n_3217: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2641,
        in1(1) => S2590,
        out1 => S2644
    );
nor_n_3218: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2641,
        in1(1) => S2590,
        out1 => S2645
    );
nand_n_3219: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2642,
        in1(1) => S2589,
        out1 => S2646
    );
nor_n_3220: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2645,
        in1(1) => S2643,
        out1 => S2648
    );
nand_n_3221: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2646,
        in1(1) => S2644,
        out1 => S2649
    );
nor_n_3222: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2649,
        in1(1) => S2588,
        out1 => S2650
    );
nand_n_3223: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2648,
        in1(1) => S2587,
        out1 => S2651
    );
nor_n_3224: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2648,
        in1(1) => S2587,
        out1 => S2652
    );
nand_n_3225: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2649,
        in1(1) => S2588,
        out1 => S2653
    );
nor_n_3226: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2652,
        in1(1) => S2650,
        out1 => S2654
    );
nand_n_3227: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2653,
        in1(1) => S2651,
        out1 => S2655
    );
nor_n_3228: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2655,
        in1(1) => S2566,
        out1 => S2656
    );
nand_n_3229: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2654,
        in1(1) => S2567,
        out1 => S2657
    );
nand_n_3230: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2655,
        in1(1) => S2566,
        out1 => S2659
    );
nand_n_3231: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2659,
        in1(1) => S2657,
        out1 => S2660
    );
notg_3232: ENTITY WORK.notg
    PORT MAP (
        in1 => S2660,
        out1 => S2661
    );
nand_n_3233: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2661,
        in1(1) => S2482,
        out1 => S2662
    );
notg_3234: ENTITY WORK.notg
    PORT MAP (
        in1 => S2662,
        out1 => S2663
    );
nand_n_3235: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2660,
        in1(1) => S2483,
        out1 => S2664
    );
nand_n_3236: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2664,
        in1(1) => S2662,
        out1 => S2665
    );
notg_3237: ENTITY WORK.notg
    PORT MAP (
        in1 => S2665,
        out1 => S2666
    );
nand_n_3238: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2666,
        in1(1) => S2552,
        out1 => S2667
    );
notg_3239: ENTITY WORK.notg
    PORT MAP (
        in1 => S2667,
        out1 => S2668
    );
nand_n_3240: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2665,
        in1(1) => S2551,
        out1 => S2670
    );
nand_n_3241: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2670,
        in1(1) => S2667,
        out1 => S2671
    );
notg_3242: ENTITY WORK.notg
    PORT MAP (
        in1 => S2671,
        out1 => S2672
    );
nand_n_3243: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2672,
        in1(1) => S2559,
        out1 => S2673
    );
nand_n_3244: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2673,
        in1(1) => S5579,
        out1 => S2674
    );
nor_n_3245: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2559,
        in1(1) => S2554,
        out1 => S2675
    );
nand_n_3246: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2675,
        in1(1) => S2671,
        out1 => S2676
    );
nand_n_3247: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2672,
        in1(1) => S2554,
        out1 => S2677
    );
nand_n_3248: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2677,
        in1(1) => S2676,
        out1 => S2678
    );
nor_n_3249: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2678,
        in1(1) => S2674,
        out1 => S2679
    );
nor_n_3250: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2679,
        in1(1) => S2564,
        out1 => S2681
    );
nand_n_3251: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2681,
        in1(1) => S2565,
        out1 => S27
    );
nor_n_3252: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S788,
        in1(1) => S5547,
        out1 => S2682
    );
nand_n_3253: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5611,
        in1(1) => new_datapath_multdivunit_outmdu1_8,
        out1 => S2683
    );
nor_n_3254: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2663,
        in1(1) => S2656,
        out1 => S2684
    );
nand_n_3255: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2662,
        in1(1) => S2657,
        out1 => S2685
    );
nor_n_3256: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2650,
        in1(1) => S2643,
        out1 => S2686
    );
nand_n_3257: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2651,
        in1(1) => S2644,
        out1 => S2687
    );
nor_n_3258: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5975,
        in1(1) => S3478,
        out1 => S2688
    );
nand_n_3259: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_0,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S2689
    );
nor_n_3260: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S202,
        in1(1) => S5957,
        out1 => S2691
    );
nand_n_3261: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S203,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S2692
    );
nor_n_3262: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2691,
        in1(1) => S2574,
        out1 => S2693
    );
nand_n_3263: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2692,
        in1(1) => S2575,
        out1 => S2694
    );
nor_n_3264: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S228,
        in1(1) => S5957,
        out1 => S2695
    );
nand_n_3265: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S229,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S2696
    );
nor_n_3266: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2692,
        in1(1) => S2575,
        out1 => S2697
    );
nand_n_3267: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2691,
        in1(1) => S2574,
        out1 => S2698
    );
nor_n_3268: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2697,
        in1(1) => S2693,
        out1 => S2699
    );
nand_n_3269: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2698,
        in1(1) => S2694,
        out1 => S2700
    );
nor_n_3270: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2700,
        in1(1) => S2689,
        out1 => S2702
    );
nand_n_3271: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2699,
        in1(1) => S2688,
        out1 => S2703
    );
nor_n_3272: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2699,
        in1(1) => S2688,
        out1 => S2704
    );
nand_n_3273: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2700,
        in1(1) => S2689,
        out1 => S2705
    );
nor_n_3274: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2704,
        in1(1) => S2702,
        out1 => S2706
    );
nand_n_3275: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2705,
        in1(1) => S2703,
        out1 => S2707
    );
nor_n_3276: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2605,
        in1(1) => S2600,
        out1 => S2708
    );
nand_n_3277: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2606,
        in1(1) => S2601,
        out1 => S2709
    );
nor_n_3278: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2708,
        in1(1) => S2707,
        out1 => S2710
    );
nand_n_3279: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2709,
        in1(1) => S2706,
        out1 => S2711
    );
nor_n_3280: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2709,
        in1(1) => S2706,
        out1 => S2713
    );
nand_n_3281: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2708,
        in1(1) => S2707,
        out1 => S2714
    );
nor_n_3282: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2713,
        in1(1) => S2710,
        out1 => S2715
    );
nand_n_3283: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2714,
        in1(1) => S2711,
        out1 => S2716
    );
nor_n_3284: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2716,
        in1(1) => S2577,
        out1 => S2717
    );
nand_n_3285: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2715,
        in1(1) => S2576,
        out1 => S2718
    );
nor_n_3286: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2715,
        in1(1) => S2576,
        out1 => S2719
    );
nand_n_3287: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2716,
        in1(1) => S2577,
        out1 => S2720
    );
nor_n_3288: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2719,
        in1(1) => S2717,
        out1 => S2721
    );
nand_n_3289: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2720,
        in1(1) => S2718,
        out1 => S2722
    );
nor_n_3290: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2637,
        in1(1) => S2630,
        out1 => S2724
    );
nand_n_3291: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2638,
        in1(1) => S2631,
        out1 => S2725
    );
nor_n_3292: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S208,
        in1(1) => S5947,
        out1 => S2726
    );
nand_n_3293: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S209,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S2727
    );
nor_n_3294: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S248,
        in1(1) => S5926,
        out1 => S2728
    );
nand_n_3295: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S249,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S2729
    );
nor_n_3296: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2728,
        in1(1) => S2598,
        out1 => S2730
    );
nand_n_3297: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2729,
        in1(1) => S2599,
        out1 => S2731
    );
nor_n_3298: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S240,
        in1(1) => S5926,
        out1 => S2732
    );
nand_n_3299: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S241,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S2733
    );
nor_n_3300: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2729,
        in1(1) => S2599,
        out1 => S2735
    );
nand_n_3301: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2728,
        in1(1) => S2598,
        out1 => S2736
    );
nor_n_3302: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2735,
        in1(1) => S2730,
        out1 => S2737
    );
nand_n_3303: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2736,
        in1(1) => S2731,
        out1 => S2738
    );
nor_n_3304: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2738,
        in1(1) => S2727,
        out1 => S2739
    );
nand_n_3305: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2737,
        in1(1) => S2726,
        out1 => S2740
    );
nor_n_3306: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2737,
        in1(1) => S2726,
        out1 => S2741
    );
nand_n_3307: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2738,
        in1(1) => S2727,
        out1 => S2742
    );
nor_n_3308: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2741,
        in1(1) => S2739,
        out1 => S2743
    );
nand_n_3309: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2742,
        in1(1) => S2740,
        out1 => S2744
    );
nor_n_3310: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2623,
        in1(1) => S2619,
        out1 => S2746
    );
nand_n_3311: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2624,
        in1(1) => S2620,
        out1 => S2747
    );
nor_n_3312: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S256,
        in1(1) => S5916,
        out1 => S2748
    );
nand_n_3313: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S2749
    );
nand_n_3314: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S2750
    );
nand_n_3315: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2750,
        in1(1) => S2618,
        out1 => S2751
    );
notg_3316: ENTITY WORK.notg
    PORT MAP (
        in1 => S2751,
        out1 => S2752
    );
nor_n_3317: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S264,
        in1(1) => S3325,
        out1 => S2753
    );
nand_n_3318: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S265,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S2754
    );
nor_n_3319: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2754,
        in1(1) => S887,
        out1 => S2755
    );
nand_n_3320: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2753,
        in1(1) => S886,
        out1 => S2757
    );
nor_n_3321: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2755,
        in1(1) => S2752,
        out1 => S2758
    );
nand_n_3322: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2757,
        in1(1) => S2751,
        out1 => S2759
    );
nor_n_3323: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2759,
        in1(1) => S2749,
        out1 => S2760
    );
nand_n_3324: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2758,
        in1(1) => S2748,
        out1 => S2761
    );
nor_n_3325: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2758,
        in1(1) => S2748,
        out1 => S2762
    );
nand_n_3326: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2759,
        in1(1) => S2749,
        out1 => S2763
    );
nor_n_3327: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2762,
        in1(1) => S2760,
        out1 => S2764
    );
nand_n_3328: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2763,
        in1(1) => S2761,
        out1 => S2765
    );
nor_n_3329: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2765,
        in1(1) => S2746,
        out1 => S2766
    );
nand_n_3330: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2764,
        in1(1) => S2747,
        out1 => S2768
    );
nor_n_3331: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2764,
        in1(1) => S2747,
        out1 => S2769
    );
nand_n_3332: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2765,
        in1(1) => S2746,
        out1 => S2770
    );
nor_n_3333: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2769,
        in1(1) => S2766,
        out1 => S2771
    );
nand_n_3334: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2770,
        in1(1) => S2768,
        out1 => S2772
    );
nor_n_3335: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2772,
        in1(1) => S2744,
        out1 => S2773
    );
nand_n_3336: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2771,
        in1(1) => S2743,
        out1 => S2774
    );
nor_n_3337: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2771,
        in1(1) => S2743,
        out1 => S2775
    );
nand_n_3338: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2772,
        in1(1) => S2744,
        out1 => S2776
    );
nor_n_3339: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2775,
        in1(1) => S2773,
        out1 => S2777
    );
nand_n_3340: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2776,
        in1(1) => S2774,
        out1 => S2779
    );
nor_n_3341: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2779,
        in1(1) => S2724,
        out1 => S2780
    );
nand_n_3342: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2777,
        in1(1) => S2725,
        out1 => S2781
    );
nor_n_3343: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2777,
        in1(1) => S2725,
        out1 => S2782
    );
nand_n_3344: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2779,
        in1(1) => S2724,
        out1 => S2783
    );
nor_n_3345: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2782,
        in1(1) => S2780,
        out1 => S2784
    );
nand_n_3346: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2783,
        in1(1) => S2781,
        out1 => S2785
    );
nor_n_3347: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2785,
        in1(1) => S2722,
        out1 => S2786
    );
nand_n_3348: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2784,
        in1(1) => S2721,
        out1 => S2787
    );
nor_n_3349: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2784,
        in1(1) => S2721,
        out1 => S2788
    );
nand_n_3350: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2785,
        in1(1) => S2722,
        out1 => S2790
    );
nor_n_3351: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2788,
        in1(1) => S2786,
        out1 => S2791
    );
nand_n_3352: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2790,
        in1(1) => S2787,
        out1 => S2792
    );
nor_n_3353: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2792,
        in1(1) => S2686,
        out1 => S2793
    );
nand_n_3354: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2791,
        in1(1) => S2687,
        out1 => S2794
    );
nor_n_3355: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2791,
        in1(1) => S2687,
        out1 => S2795
    );
nand_n_3356: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2792,
        in1(1) => S2686,
        out1 => S2796
    );
nor_n_3357: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2795,
        in1(1) => S2793,
        out1 => S2797
    );
nand_n_3358: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2796,
        in1(1) => S2794,
        out1 => S2798
    );
nor_n_3359: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2798,
        in1(1) => S2586,
        out1 => S2799
    );
nand_n_3360: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2797,
        in1(1) => S2585,
        out1 => S2801
    );
nor_n_3361: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2797,
        in1(1) => S2585,
        out1 => S2802
    );
nand_n_3362: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2798,
        in1(1) => S2586,
        out1 => S2803
    );
nor_n_3363: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2802,
        in1(1) => S2799,
        out1 => S2804
    );
nand_n_3364: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2803,
        in1(1) => S2801,
        out1 => S2805
    );
nand_n_3365: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2805,
        in1(1) => S2684,
        out1 => S2806
    );
nor_n_3366: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2805,
        in1(1) => S2684,
        out1 => S2807
    );
nand_n_3367: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2804,
        in1(1) => S2685,
        out1 => S2808
    );
nand_n_3368: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2808,
        in1(1) => S2806,
        out1 => S2809
    );
notg_3369: ENTITY WORK.notg
    PORT MAP (
        in1 => S2809,
        out1 => S2810
    );
nand_n_3370: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2810,
        in1(1) => S2668,
        out1 => S2812
    );
notg_3371: ENTITY WORK.notg
    PORT MAP (
        in1 => S2812,
        out1 => S2813
    );
nand_n_3372: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2809,
        in1(1) => S2667,
        out1 => S2814
    );
nand_n_3373: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2814,
        in1(1) => S2812,
        out1 => S2815
    );
nor_n_3374: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2815,
        in1(1) => S2677,
        out1 => S2816
    );
notg_3375: ENTITY WORK.notg
    PORT MAP (
        in1 => S2816,
        out1 => S2817
    );
nand_n_3376: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2815,
        in1(1) => S2677,
        out1 => S2818
    );
nand_n_3377: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2818,
        in1(1) => S2817,
        out1 => S2819
    );
nor_n_3378: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2819,
        in1(1) => S2673,
        out1 => S2820
    );
nand_n_3379: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2819,
        in1(1) => S2673,
        out1 => S2821
    );
nand_n_3380: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2821,
        in1(1) => S5579,
        out1 => S2823
    );
nor_n_3381: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2823,
        in1(1) => S2820,
        out1 => S2824
    );
nor_n_3382: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2824,
        in1(1) => S2682,
        out1 => S2825
    );
nand_n_3383: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2825,
        in1(1) => S2683,
        out1 => S28
    );
nor_n_3384: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S664,
        in1(1) => S5547,
        out1 => S2826
    );
nand_n_3385: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5611,
        in1(1) => new_datapath_multdivunit_outmdu1_9,
        out1 => S2827
    );
nor_n_3386: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2820,
        in1(1) => S2816,
        out1 => S2828
    );
nor_n_3387: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2799,
        in1(1) => S2793,
        out1 => S2829
    );
nand_n_3388: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2801,
        in1(1) => S2794,
        out1 => S2830
    );
nor_n_3389: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5975,
        in1(1) => S3467,
        out1 => S2831
    );
nand_n_3390: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_0,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S2833
    );
nor_n_3391: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2717,
        in1(1) => S2710,
        out1 => S2834
    );
nand_n_3392: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2718,
        in1(1) => S2711,
        out1 => S2835
    );
nor_n_3393: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2834,
        in1(1) => S2833,
        out1 => S2836
    );
nand_n_3394: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2835,
        in1(1) => S2831,
        out1 => S2837
    );
nor_n_3395: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2835,
        in1(1) => S2831,
        out1 => S2838
    );
nand_n_3396: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2834,
        in1(1) => S2833,
        out1 => S2839
    );
nor_n_3397: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2838,
        in1(1) => S2836,
        out1 => S2840
    );
nand_n_3398: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2839,
        in1(1) => S2837,
        out1 => S2841
    );
nor_n_3399: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2786,
        in1(1) => S2780,
        out1 => S2842
    );
nand_n_3400: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2787,
        in1(1) => S2781,
        out1 => S2844
    );
nor_n_3401: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2702,
        in1(1) => S2697,
        out1 => S2845
    );
nand_n_3402: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2703,
        in1(1) => S2698,
        out1 => S2846
    );
nor_n_3403: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5966,
        in1(1) => S3478,
        out1 => S2847
    );
nand_n_3404: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_1,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S2848
    );
nor_n_3405: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S202,
        in1(1) => S5947,
        out1 => S2849
    );
nand_n_3406: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S203,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S2850
    );
nor_n_3407: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2849,
        in1(1) => S2695,
        out1 => S2851
    );
nand_n_3408: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2850,
        in1(1) => S2696,
        out1 => S2852
    );
nor_n_3409: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S228,
        in1(1) => S5947,
        out1 => S2853
    );
nand_n_3410: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S229,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S2855
    );
nor_n_3411: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2850,
        in1(1) => S2696,
        out1 => S2856
    );
nand_n_3412: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2849,
        in1(1) => S2695,
        out1 => S2857
    );
nor_n_3413: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2856,
        in1(1) => S2851,
        out1 => S2858
    );
nand_n_3414: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2857,
        in1(1) => S2852,
        out1 => S2859
    );
nor_n_3415: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2859,
        in1(1) => S2848,
        out1 => S2860
    );
nand_n_3416: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2858,
        in1(1) => S2847,
        out1 => S2861
    );
nor_n_3417: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2858,
        in1(1) => S2847,
        out1 => S2862
    );
nand_n_3418: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2859,
        in1(1) => S2848,
        out1 => S2863
    );
nor_n_3419: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2862,
        in1(1) => S2860,
        out1 => S2864
    );
nand_n_3420: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2863,
        in1(1) => S2861,
        out1 => S2866
    );
nor_n_3421: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2739,
        in1(1) => S2735,
        out1 => S2867
    );
nand_n_3422: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2740,
        in1(1) => S2736,
        out1 => S2868
    );
nor_n_3423: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2867,
        in1(1) => S2866,
        out1 => S2869
    );
nand_n_3424: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2868,
        in1(1) => S2864,
        out1 => S2870
    );
nor_n_3425: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2868,
        in1(1) => S2864,
        out1 => S2871
    );
nand_n_3426: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2867,
        in1(1) => S2866,
        out1 => S2872
    );
nor_n_3427: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2871,
        in1(1) => S2869,
        out1 => S2873
    );
nand_n_3428: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2872,
        in1(1) => S2870,
        out1 => S2874
    );
nor_n_3429: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2873,
        in1(1) => S2846,
        out1 => S2875
    );
nand_n_3430: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2874,
        in1(1) => S2845,
        out1 => S2877
    );
nor_n_3431: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2874,
        in1(1) => S2845,
        out1 => S2878
    );
nand_n_3432: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2873,
        in1(1) => S2846,
        out1 => S2879
    );
nor_n_3433: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2878,
        in1(1) => S2875,
        out1 => S2880
    );
nand_n_3434: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2879,
        in1(1) => S2877,
        out1 => S2881
    );
nor_n_3435: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2773,
        in1(1) => S2766,
        out1 => S2882
    );
nand_n_3436: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2774,
        in1(1) => S2768,
        out1 => S2883
    );
nor_n_3437: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S208,
        in1(1) => S5936,
        out1 => S2884
    );
nand_n_3438: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S209,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S2885
    );
nor_n_3439: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S248,
        in1(1) => S5916,
        out1 => S2886
    );
nand_n_3440: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S249,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S2888
    );
nor_n_3441: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2886,
        in1(1) => S2732,
        out1 => S2889
    );
nand_n_3442: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2888,
        in1(1) => S2733,
        out1 => S2890
    );
nor_n_3443: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S240,
        in1(1) => S5916,
        out1 => S2891
    );
nand_n_3444: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S241,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S2892
    );
nor_n_3445: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2888,
        in1(1) => S2733,
        out1 => S2893
    );
nand_n_3446: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2886,
        in1(1) => S2732,
        out1 => S2894
    );
nor_n_3447: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2893,
        in1(1) => S2889,
        out1 => S2895
    );
nand_n_3448: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2894,
        in1(1) => S2890,
        out1 => S2896
    );
nor_n_3449: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2896,
        in1(1) => S2885,
        out1 => S2897
    );
nand_n_3450: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2895,
        in1(1) => S2884,
        out1 => S2899
    );
nor_n_3451: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2895,
        in1(1) => S2884,
        out1 => S2900
    );
nand_n_3452: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2896,
        in1(1) => S2885,
        out1 => S2901
    );
nor_n_3453: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2900,
        in1(1) => S2897,
        out1 => S2902
    );
nand_n_3454: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2901,
        in1(1) => S2899,
        out1 => S2903
    );
nor_n_3455: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2760,
        in1(1) => S2755,
        out1 => S2904
    );
nand_n_3456: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2761,
        in1(1) => S2757,
        out1 => S2905
    );
nor_n_3457: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S256,
        in1(1) => S5907,
        out1 => S2906
    );
nand_n_3458: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S2907
    );
nor_n_3459: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2753,
        in1(1) => S736,
        out1 => S2908
    );
nand_n_3460: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2754,
        in1(1) => S737,
        out1 => S2910
    );
nand_n_3461: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S265,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S2911
    );
nor_n_3462: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2754,
        in1(1) => S737,
        out1 => S2912
    );
nand_n_3463: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2753,
        in1(1) => S736,
        out1 => S2913
    );
nor_n_3464: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2912,
        in1(1) => S2908,
        out1 => S2914
    );
nand_n_3465: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2913,
        in1(1) => S2910,
        out1 => S2915
    );
nor_n_3466: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2915,
        in1(1) => S2907,
        out1 => S2916
    );
nand_n_3467: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2914,
        in1(1) => S2906,
        out1 => S2917
    );
nor_n_3468: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2914,
        in1(1) => S2906,
        out1 => S2918
    );
nand_n_3469: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2915,
        in1(1) => S2907,
        out1 => S2919
    );
nor_n_3470: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2918,
        in1(1) => S2916,
        out1 => S2921
    );
nand_n_3471: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2919,
        in1(1) => S2917,
        out1 => S2922
    );
nor_n_3472: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2922,
        in1(1) => S2904,
        out1 => S2923
    );
nand_n_3473: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2921,
        in1(1) => S2905,
        out1 => S2924
    );
nor_n_3474: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2921,
        in1(1) => S2905,
        out1 => S2925
    );
nand_n_3475: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2922,
        in1(1) => S2904,
        out1 => S2926
    );
nor_n_3476: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2925,
        in1(1) => S2923,
        out1 => S2927
    );
nand_n_3477: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2926,
        in1(1) => S2924,
        out1 => S2928
    );
nor_n_3478: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2928,
        in1(1) => S2903,
        out1 => S2929
    );
nand_n_3479: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2927,
        in1(1) => S2902,
        out1 => S2930
    );
nor_n_3480: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2927,
        in1(1) => S2902,
        out1 => S2932
    );
nand_n_3481: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2928,
        in1(1) => S2903,
        out1 => S2933
    );
nor_n_3482: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2932,
        in1(1) => S2929,
        out1 => S2934
    );
nand_n_3483: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2933,
        in1(1) => S2930,
        out1 => S2935
    );
nor_n_3484: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2935,
        in1(1) => S2882,
        out1 => S2936
    );
nand_n_3485: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2934,
        in1(1) => S2883,
        out1 => S2937
    );
nor_n_3486: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2934,
        in1(1) => S2883,
        out1 => S2938
    );
nand_n_3487: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2935,
        in1(1) => S2882,
        out1 => S2939
    );
nor_n_3488: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2938,
        in1(1) => S2936,
        out1 => S2940
    );
nand_n_3489: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2939,
        in1(1) => S2937,
        out1 => S2941
    );
nor_n_3490: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2941,
        in1(1) => S2881,
        out1 => S2943
    );
nand_n_3491: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2940,
        in1(1) => S2880,
        out1 => S2944
    );
nor_n_3492: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2940,
        in1(1) => S2880,
        out1 => S2945
    );
nand_n_3493: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2941,
        in1(1) => S2881,
        out1 => S2946
    );
nor_n_3494: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2945,
        in1(1) => S2943,
        out1 => S2947
    );
nand_n_3495: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2946,
        in1(1) => S2944,
        out1 => S2948
    );
nor_n_3496: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2948,
        in1(1) => S2842,
        out1 => S2949
    );
nand_n_3497: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2947,
        in1(1) => S2844,
        out1 => S2950
    );
nor_n_3498: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2947,
        in1(1) => S2844,
        out1 => S2951
    );
nand_n_3499: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2948,
        in1(1) => S2842,
        out1 => S2952
    );
nor_n_3500: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2951,
        in1(1) => S2949,
        out1 => S2954
    );
nand_n_3501: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2952,
        in1(1) => S2950,
        out1 => S2955
    );
nor_n_3502: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2955,
        in1(1) => S2841,
        out1 => S2956
    );
nand_n_3503: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2954,
        in1(1) => S2840,
        out1 => S2957
    );
nor_n_3504: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2954,
        in1(1) => S2840,
        out1 => S2958
    );
nand_n_3505: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2955,
        in1(1) => S2841,
        out1 => S2959
    );
nor_n_3506: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2958,
        in1(1) => S2956,
        out1 => S2960
    );
nand_n_3507: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2959,
        in1(1) => S2957,
        out1 => S2961
    );
nor_n_3508: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2960,
        in1(1) => S2830,
        out1 => S2962
    );
nand_n_3509: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2961,
        in1(1) => S2829,
        out1 => S2963
    );
nor_n_3510: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2961,
        in1(1) => S2829,
        out1 => S2965
    );
notg_3511: ENTITY WORK.notg
    PORT MAP (
        in1 => S2965,
        out1 => S2966
    );
nor_n_3512: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2965,
        in1(1) => S2962,
        out1 => S2967
    );
nand_n_3513: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2966,
        in1(1) => S2963,
        out1 => S2968
    );
nor_n_3514: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2968,
        in1(1) => S2808,
        out1 => S2969
    );
nand_n_3515: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2967,
        in1(1) => S2807,
        out1 => S2970
    );
nor_n_3516: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2967,
        in1(1) => S2807,
        out1 => S2971
    );
nand_n_3517: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2968,
        in1(1) => S2808,
        out1 => S2972
    );
nor_n_3518: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2971,
        in1(1) => S2969,
        out1 => S2973
    );
nand_n_3519: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2972,
        in1(1) => S2970,
        out1 => S2974
    );
nand_n_3520: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2973,
        in1(1) => S2813,
        out1 => S2976
    );
nand_n_3521: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2974,
        in1(1) => S2812,
        out1 => S2977
    );
nand_n_3522: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2977,
        in1(1) => S2976,
        out1 => S2978
    );
nor_n_3523: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2978,
        in1(1) => S2828,
        out1 => S2979
    );
notg_3524: ENTITY WORK.notg
    PORT MAP (
        in1 => S2979,
        out1 => S2980
    );
nand_n_3525: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2978,
        in1(1) => S2828,
        out1 => S2981
    );
nand_n_3526: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2981,
        in1(1) => S5579,
        out1 => S2982
    );
nor_n_3527: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2982,
        in1(1) => S2979,
        out1 => S2983
    );
nor_n_3528: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2983,
        in1(1) => S2826,
        out1 => S2984
    );
nand_n_3529: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2984,
        in1(1) => S2827,
        out1 => S29
    );
nor_n_3530: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S557,
        in1(1) => S5547,
        out1 => S2986
    );
nand_n_3531: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5611,
        in1(1) => new_datapath_multdivunit_outmdu1_10,
        out1 => S2987
    );
nand_n_3532: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2980,
        in1(1) => S2976,
        out1 => S2988
    );
nor_n_3533: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2956,
        in1(1) => S2949,
        out1 => S2989
    );
nand_n_3534: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2957,
        in1(1) => S2950,
        out1 => S2990
    );
nand_n_3535: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_0,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S2991
    );
nand_n_3536: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_1,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S2992
    );
nand_n_3537: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2992,
        in1(1) => S2991,
        out1 => S2993
    );
notg_3538: ENTITY WORK.notg
    PORT MAP (
        in1 => S2993,
        out1 => S2994
    );
nor_n_3539: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5966,
        in1(1) => S3456,
        out1 => S2995
    );
nand_n_3540: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_1,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S2997
    );
nor_n_3541: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2997,
        in1(1) => S2833,
        out1 => S2998
    );
nand_n_3542: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2995,
        in1(1) => S2831,
        out1 => S2999
    );
nor_n_3543: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2998,
        in1(1) => S2994,
        out1 => S3000
    );
nand_n_3544: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2999,
        in1(1) => S2993,
        out1 => S3001
    );
nor_n_3545: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2878,
        in1(1) => S2869,
        out1 => S3002
    );
nand_n_3546: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2879,
        in1(1) => S2870,
        out1 => S3003
    );
nor_n_3547: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3003,
        in1(1) => S3000,
        out1 => S3004
    );
nand_n_3548: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3002,
        in1(1) => S3001,
        out1 => S3005
    );
nor_n_3549: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3002,
        in1(1) => S3001,
        out1 => S3006
    );
nand_n_3550: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3003,
        in1(1) => S3000,
        out1 => S3008
    );
nor_n_3551: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3006,
        in1(1) => S3004,
        out1 => S3009
    );
nand_n_3552: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3008,
        in1(1) => S3005,
        out1 => S3010
    );
nor_n_3553: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2943,
        in1(1) => S2936,
        out1 => S3011
    );
nand_n_3554: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2944,
        in1(1) => S2937,
        out1 => S3012
    );
nor_n_3555: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2860,
        in1(1) => S2856,
        out1 => S3013
    );
nand_n_3556: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2861,
        in1(1) => S2857,
        out1 => S3014
    );
nor_n_3557: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5957,
        in1(1) => S3478,
        out1 => S3015
    );
nand_n_3558: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_2,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S3016
    );
nor_n_3559: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S202,
        in1(1) => S5936,
        out1 => S3017
    );
nand_n_3560: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S203,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S3019
    );
nor_n_3561: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3017,
        in1(1) => S2853,
        out1 => S3020
    );
nand_n_3562: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3019,
        in1(1) => S2855,
        out1 => S3021
    );
nor_n_3563: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S228,
        in1(1) => S5936,
        out1 => S3022
    );
nand_n_3564: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S229,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S3023
    );
nor_n_3565: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3019,
        in1(1) => S2855,
        out1 => S3024
    );
nand_n_3566: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3017,
        in1(1) => S2853,
        out1 => S3025
    );
nor_n_3567: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3024,
        in1(1) => S3020,
        out1 => S3026
    );
nand_n_3568: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3025,
        in1(1) => S3021,
        out1 => S3027
    );
nor_n_3569: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3027,
        in1(1) => S3016,
        out1 => S3028
    );
nand_n_3570: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3026,
        in1(1) => S3015,
        out1 => S3030
    );
nor_n_3571: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3026,
        in1(1) => S3015,
        out1 => S3031
    );
nand_n_3572: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3027,
        in1(1) => S3016,
        out1 => S3032
    );
nor_n_3573: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3031,
        in1(1) => S3028,
        out1 => S3033
    );
nand_n_3574: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3032,
        in1(1) => S3030,
        out1 => S3034
    );
nor_n_3575: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2897,
        in1(1) => S2893,
        out1 => S3035
    );
nand_n_3576: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2899,
        in1(1) => S2894,
        out1 => S3036
    );
nor_n_3577: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3035,
        in1(1) => S3034,
        out1 => S3037
    );
nand_n_3578: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3036,
        in1(1) => S3033,
        out1 => S3038
    );
nor_n_3579: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3036,
        in1(1) => S3033,
        out1 => S3039
    );
nand_n_3580: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3035,
        in1(1) => S3034,
        out1 => S3041
    );
nor_n_3581: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3039,
        in1(1) => S3037,
        out1 => S3042
    );
nand_n_3582: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3041,
        in1(1) => S3038,
        out1 => S3043
    );
nor_n_3583: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3042,
        in1(1) => S3014,
        out1 => S3044
    );
nand_n_3584: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3043,
        in1(1) => S3013,
        out1 => S3045
    );
nor_n_3585: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3043,
        in1(1) => S3013,
        out1 => S3046
    );
nand_n_3586: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3042,
        in1(1) => S3014,
        out1 => S3047
    );
nor_n_3587: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3046,
        in1(1) => S3044,
        out1 => S3048
    );
nand_n_3588: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3047,
        in1(1) => S3045,
        out1 => S3049
    );
nor_n_3589: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2929,
        in1(1) => S2923,
        out1 => S3050
    );
nand_n_3590: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2930,
        in1(1) => S2924,
        out1 => S3052
    );
nor_n_3591: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S208,
        in1(1) => S5926,
        out1 => S3053
    );
nand_n_3592: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S209,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S3054
    );
nor_n_3593: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S248,
        in1(1) => S5907,
        out1 => S3055
    );
nand_n_3594: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S249,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S3056
    );
nor_n_3595: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3055,
        in1(1) => S2891,
        out1 => S3057
    );
nand_n_3596: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3056,
        in1(1) => S2892,
        out1 => S3058
    );
nor_n_3597: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S240,
        in1(1) => S5907,
        out1 => S3059
    );
nand_n_3598: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S241,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S3060
    );
nor_n_3599: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3056,
        in1(1) => S2892,
        out1 => S3061
    );
nand_n_3600: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3055,
        in1(1) => S2891,
        out1 => S3063
    );
nor_n_3601: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3061,
        in1(1) => S3057,
        out1 => S3064
    );
nand_n_3602: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3063,
        in1(1) => S3058,
        out1 => S3065
    );
nor_n_3603: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3065,
        in1(1) => S3054,
        out1 => S3066
    );
nand_n_3604: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3064,
        in1(1) => S3053,
        out1 => S3067
    );
nor_n_3605: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3064,
        in1(1) => S3053,
        out1 => S3068
    );
nand_n_3606: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3065,
        in1(1) => S3054,
        out1 => S3069
    );
nor_n_3607: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3068,
        in1(1) => S3066,
        out1 => S3070
    );
nand_n_3608: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3069,
        in1(1) => S3067,
        out1 => S3071
    );
nor_n_3609: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S2916,
        in1(1) => S2912,
        out1 => S3072
    );
nand_n_3610: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S2917,
        in1(1) => S2913,
        out1 => S3074
    );
nand_n_3611: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S3075
    );
notg_3612: ENTITY WORK.notg
    PORT MAP (
        in1 => S3075,
        out1 => S3076
    );
nand_n_3613: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S3077
    );
nand_n_3614: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3077,
        in1(1) => S2911,
        out1 => S3078
    );
nor_n_3615: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S264,
        in1(1) => S3346,
        out1 => S3079
    );
nand_n_3616: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S265,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S3080
    );
nor_n_3617: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3080,
        in1(1) => S737,
        out1 => S3081
    );
nand_n_3618: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3079,
        in1(1) => S736,
        out1 => S3082
    );
nand_n_3619: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3082,
        in1(1) => S3078,
        out1 => S3083
    );
notg_3620: ENTITY WORK.notg
    PORT MAP (
        in1 => S3083,
        out1 => S3085
    );
nor_n_3621: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3083,
        in1(1) => S3075,
        out1 => S3086
    );
nand_n_3622: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3085,
        in1(1) => S3076,
        out1 => S3087
    );
nand_n_3623: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3083,
        in1(1) => S3075,
        out1 => S3088
    );
notg_3624: ENTITY WORK.notg
    PORT MAP (
        in1 => S3088,
        out1 => S3089
    );
nor_n_3625: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3089,
        in1(1) => S3086,
        out1 => S3090
    );
nand_n_3626: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3088,
        in1(1) => S3087,
        out1 => S3091
    );
nor_n_3627: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3091,
        in1(1) => S3072,
        out1 => S3092
    );
nand_n_3628: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3090,
        in1(1) => S3074,
        out1 => S3093
    );
nor_n_3629: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3090,
        in1(1) => S3074,
        out1 => S3094
    );
nand_n_3630: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3091,
        in1(1) => S3072,
        out1 => S3096
    );
nor_n_3631: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3094,
        in1(1) => S3092,
        out1 => S3097
    );
nand_n_3632: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3096,
        in1(1) => S3093,
        out1 => S3098
    );
nor_n_3633: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3098,
        in1(1) => S3071,
        out1 => S3099
    );
nand_n_3634: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3097,
        in1(1) => S3070,
        out1 => S3100
    );
nor_n_3635: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3097,
        in1(1) => S3070,
        out1 => S3101
    );
nand_n_3636: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3098,
        in1(1) => S3071,
        out1 => S3102
    );
nor_n_3637: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3101,
        in1(1) => S3099,
        out1 => S3103
    );
nand_n_3638: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3102,
        in1(1) => S3100,
        out1 => S3104
    );
nor_n_3639: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3104,
        in1(1) => S3050,
        out1 => S3105
    );
nand_n_3640: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3103,
        in1(1) => S3052,
        out1 => S3107
    );
nor_n_3641: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3103,
        in1(1) => S3052,
        out1 => S3108
    );
nand_n_3642: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3104,
        in1(1) => S3050,
        out1 => S3109
    );
nor_n_3643: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3108,
        in1(1) => S3105,
        out1 => S3110
    );
nand_n_3644: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3109,
        in1(1) => S3107,
        out1 => S3111
    );
nor_n_3645: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3111,
        in1(1) => S3049,
        out1 => S3112
    );
nand_n_3646: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3110,
        in1(1) => S3048,
        out1 => S3113
    );
nor_n_3647: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3110,
        in1(1) => S3048,
        out1 => S3114
    );
nand_n_3648: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3111,
        in1(1) => S3049,
        out1 => S3115
    );
nor_n_3649: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3114,
        in1(1) => S3112,
        out1 => S3116
    );
nand_n_3650: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3115,
        in1(1) => S3113,
        out1 => S3118
    );
nor_n_3651: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3118,
        in1(1) => S3011,
        out1 => S3119
    );
nand_n_3652: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3116,
        in1(1) => S3012,
        out1 => S3120
    );
nor_n_3653: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3116,
        in1(1) => S3012,
        out1 => S3121
    );
nand_n_3654: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3118,
        in1(1) => S3011,
        out1 => S3122
    );
nor_n_3655: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3121,
        in1(1) => S3119,
        out1 => S3123
    );
nand_n_3656: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3122,
        in1(1) => S3120,
        out1 => S3124
    );
nor_n_3657: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3124,
        in1(1) => S3010,
        out1 => S3125
    );
nand_n_3658: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3123,
        in1(1) => S3009,
        out1 => S3126
    );
nor_n_3659: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3123,
        in1(1) => S3009,
        out1 => S3127
    );
nand_n_3660: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3124,
        in1(1) => S3010,
        out1 => S3129
    );
nor_n_3661: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3127,
        in1(1) => S3125,
        out1 => S3130
    );
nand_n_3662: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3129,
        in1(1) => S3126,
        out1 => S3131
    );
nor_n_3663: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3131,
        in1(1) => S2989,
        out1 => S3132
    );
nand_n_3664: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3130,
        in1(1) => S2990,
        out1 => S3133
    );
nor_n_3665: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3130,
        in1(1) => S2990,
        out1 => S3134
    );
nand_n_3666: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3131,
        in1(1) => S2989,
        out1 => S3135
    );
nor_n_3667: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3134,
        in1(1) => S3132,
        out1 => S3136
    );
nand_n_3668: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3135,
        in1(1) => S3133,
        out1 => S3137
    );
nor_n_3669: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3137,
        in1(1) => S2837,
        out1 => S3138
    );
nor_n_3670: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3136,
        in1(1) => S2836,
        out1 => S3140
    );
nor_n_3671: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3140,
        in1(1) => S3138,
        out1 => S3141
    );
nand_n_3672: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3141,
        in1(1) => S2965,
        out1 => S3142
    );
notg_3673: ENTITY WORK.notg
    PORT MAP (
        in1 => S3142,
        out1 => S3143
    );
nor_n_3674: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3141,
        in1(1) => S2965,
        out1 => S3144
    );
notg_3675: ENTITY WORK.notg
    PORT MAP (
        in1 => S3144,
        out1 => S3145
    );
nor_n_3676: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3144,
        in1(1) => S3143,
        out1 => S3146
    );
nand_n_3677: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3145,
        in1(1) => S3142,
        out1 => S3147
    );
nor_n_3678: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3147,
        in1(1) => S2970,
        out1 => S3148
    );
nor_n_3679: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3146,
        in1(1) => S2969,
        out1 => S3149
    );
nor_n_3680: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3149,
        in1(1) => S3148,
        out1 => S3151
    );
nand_n_3681: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3151,
        in1(1) => S2988,
        out1 => S3152
    );
notg_3682: ENTITY WORK.notg
    PORT MAP (
        in1 => S3152,
        out1 => S3153
    );
nor_n_3683: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3151,
        in1(1) => S2988,
        out1 => S3154
    );
nand_n_3684: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3152,
        in1(1) => S5579,
        out1 => S3155
    );
nor_n_3685: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3155,
        in1(1) => S3154,
        out1 => S3156
    );
nor_n_3686: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3156,
        in1(1) => S2986,
        out1 => S3157
    );
nand_n_3687: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3157,
        in1(1) => S2987,
        out1 => S30
    );
nor_n_3688: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S461,
        in1(1) => S5547,
        out1 => S3158
    );
nand_n_3689: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5611,
        in1(1) => new_datapath_multdivunit_outmdu1_11,
        out1 => S3159
    );
nor_n_3690: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3153,
        in1(1) => S3148,
        out1 => S3161
    );
nor_n_3691: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3138,
        in1(1) => S3132,
        out1 => S3162
    );
notg_3692: ENTITY WORK.notg
    PORT MAP (
        in1 => S3162,
        out1 => S3163
    );
nor_n_3693: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3125,
        in1(1) => S3119,
        out1 => S3164
    );
nand_n_3694: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3126,
        in1(1) => S3120,
        out1 => S3165
    );
nand_n_3695: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_0,
        in1(1) => new_datapath_multdivunit_1697_B_11,
        out1 => S3166
    );
notg_3696: ENTITY WORK.notg
    PORT MAP (
        in1 => S3166,
        out1 => S3167
    );
nor_n_3697: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5957,
        in1(1) => S3467,
        out1 => S3168
    );
nand_n_3698: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_2,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S3169
    );
nand_n_3699: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3169,
        in1(1) => S2997,
        out1 => S3170
    );
nand_n_3700: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_2,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S3172
    );
nor_n_3701: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3169,
        in1(1) => S2997,
        out1 => S3173
    );
nand_n_3702: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3168,
        in1(1) => S2995,
        out1 => S3174
    );
nand_n_3703: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3174,
        in1(1) => S3170,
        out1 => S3175
    );
notg_3704: ENTITY WORK.notg
    PORT MAP (
        in1 => S3175,
        out1 => S3176
    );
nor_n_3705: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3175,
        in1(1) => S3166,
        out1 => S3177
    );
nand_n_3706: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3176,
        in1(1) => S3167,
        out1 => S3178
    );
nand_n_3707: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3175,
        in1(1) => S3166,
        out1 => S3179
    );
notg_3708: ENTITY WORK.notg
    PORT MAP (
        in1 => S3179,
        out1 => S3180
    );
nor_n_3709: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3180,
        in1(1) => S3177,
        out1 => S3181
    );
nand_n_3710: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3179,
        in1(1) => S3178,
        out1 => S3183
    );
nor_n_3711: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3183,
        in1(1) => S2999,
        out1 => S3184
    );
nand_n_3712: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3181,
        in1(1) => S2998,
        out1 => S3185
    );
nor_n_3713: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3181,
        in1(1) => S2998,
        out1 => S3186
    );
nand_n_3714: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3183,
        in1(1) => S2999,
        out1 => S3187
    );
nor_n_3715: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3186,
        in1(1) => S3184,
        out1 => S3188
    );
nand_n_3716: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3187,
        in1(1) => S3185,
        out1 => S3189
    );
nor_n_3717: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3046,
        in1(1) => S3037,
        out1 => S3190
    );
nand_n_3718: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3047,
        in1(1) => S3038,
        out1 => S3191
    );
nor_n_3719: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3191,
        in1(1) => S3188,
        out1 => S3192
    );
nand_n_3720: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3190,
        in1(1) => S3189,
        out1 => S3194
    );
nor_n_3721: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3190,
        in1(1) => S3189,
        out1 => S3195
    );
nand_n_3722: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3191,
        in1(1) => S3188,
        out1 => S3196
    );
nor_n_3723: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3195,
        in1(1) => S3192,
        out1 => S3197
    );
nand_n_3724: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3196,
        in1(1) => S3194,
        out1 => S3198
    );
nor_n_3725: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3112,
        in1(1) => S3105,
        out1 => S3199
    );
nand_n_3726: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3113,
        in1(1) => S3107,
        out1 => S3200
    );
nor_n_3727: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3028,
        in1(1) => S3024,
        out1 => S3201
    );
nand_n_3728: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3030,
        in1(1) => S3025,
        out1 => S3202
    );
nor_n_3729: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5947,
        in1(1) => S3478,
        out1 => S3203
    );
nand_n_3730: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_3,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S3205
    );
nor_n_3731: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S202,
        in1(1) => S5926,
        out1 => S3206
    );
nand_n_3732: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S203,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S3207
    );
nor_n_3733: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3206,
        in1(1) => S3022,
        out1 => S3208
    );
nand_n_3734: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3207,
        in1(1) => S3023,
        out1 => S3209
    );
nor_n_3735: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S228,
        in1(1) => S5926,
        out1 => S3210
    );
nand_n_3736: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S229,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S3211
    );
nor_n_3737: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3207,
        in1(1) => S3023,
        out1 => S3212
    );
nand_n_3738: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3206,
        in1(1) => S3022,
        out1 => S3213
    );
nor_n_3739: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3212,
        in1(1) => S3208,
        out1 => S3214
    );
nand_n_3740: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3213,
        in1(1) => S3209,
        out1 => S3216
    );
nor_n_3741: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3216,
        in1(1) => S3205,
        out1 => S3217
    );
nand_n_3742: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3214,
        in1(1) => S3203,
        out1 => S3218
    );
nor_n_3743: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3214,
        in1(1) => S3203,
        out1 => S3219
    );
nand_n_3744: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3216,
        in1(1) => S3205,
        out1 => S3220
    );
nor_n_3745: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3219,
        in1(1) => S3217,
        out1 => S3221
    );
nand_n_3746: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3220,
        in1(1) => S3218,
        out1 => S3222
    );
nor_n_3747: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3066,
        in1(1) => S3061,
        out1 => S3223
    );
nand_n_3748: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3067,
        in1(1) => S3063,
        out1 => S3224
    );
nor_n_3749: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3223,
        in1(1) => S3222,
        out1 => S3225
    );
nand_n_3750: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3224,
        in1(1) => S3221,
        out1 => S3227
    );
nor_n_3751: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3224,
        in1(1) => S3221,
        out1 => S3228
    );
nand_n_3752: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3223,
        in1(1) => S3222,
        out1 => S3229
    );
nor_n_3753: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3228,
        in1(1) => S3225,
        out1 => S3230
    );
nand_n_3754: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3229,
        in1(1) => S3227,
        out1 => S3231
    );
nor_n_3755: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3230,
        in1(1) => S3202,
        out1 => S3232
    );
nand_n_3756: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3231,
        in1(1) => S3201,
        out1 => S3233
    );
nor_n_3757: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3231,
        in1(1) => S3201,
        out1 => S3234
    );
nand_n_3758: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3230,
        in1(1) => S3202,
        out1 => S3235
    );
nor_n_3759: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3234,
        in1(1) => S3232,
        out1 => S3236
    );
nand_n_3760: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3235,
        in1(1) => S3233,
        out1 => S3238
    );
nor_n_3761: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3099,
        in1(1) => S3092,
        out1 => S3239
    );
nand_n_3762: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3100,
        in1(1) => S3093,
        out1 => S3240
    );
nor_n_3763: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S208,
        in1(1) => S5916,
        out1 => S3241
    );
nand_n_3764: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S209,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S3242
    );
nor_n_3765: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S248,
        in1(1) => S3325,
        out1 => S3243
    );
nand_n_3766: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S249,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S3244
    );
nor_n_3767: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3243,
        in1(1) => S3059,
        out1 => S3245
    );
nand_n_3768: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3244,
        in1(1) => S3060,
        out1 => S3246
    );
nand_n_3769: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S241,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S3247
    );
nor_n_3770: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3244,
        in1(1) => S3060,
        out1 => S3249
    );
nand_n_3771: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3243,
        in1(1) => S3059,
        out1 => S3250
    );
nor_n_3772: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3249,
        in1(1) => S3245,
        out1 => S3251
    );
nand_n_3773: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3250,
        in1(1) => S3246,
        out1 => S3252
    );
nor_n_3774: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3252,
        in1(1) => S3242,
        out1 => S3253
    );
nand_n_3775: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3251,
        in1(1) => S3241,
        out1 => S3254
    );
nor_n_3776: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3251,
        in1(1) => S3241,
        out1 => S3255
    );
nand_n_3777: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3252,
        in1(1) => S3242,
        out1 => S3256
    );
nor_n_3778: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3255,
        in1(1) => S3253,
        out1 => S3257
    );
nand_n_3779: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3256,
        in1(1) => S3254,
        out1 => S3258
    );
nor_n_3780: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3086,
        in1(1) => S3081,
        out1 => S3260
    );
nand_n_3781: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3087,
        in1(1) => S3082,
        out1 => S3261
    );
nor_n_3782: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S256,
        in1(1) => S3336,
        out1 => S3262
    );
nand_n_3783: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S3263
    );
nor_n_3784: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3079,
        in1(1) => S511,
        out1 => S3264
    );
nand_n_3785: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3080,
        in1(1) => S512,
        out1 => S3265
    );
nand_n_3786: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S265,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S3266
    );
nor_n_3787: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3080,
        in1(1) => S512,
        out1 => S3267
    );
nand_n_3788: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3079,
        in1(1) => S511,
        out1 => S3268
    );
nor_n_3789: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3267,
        in1(1) => S3264,
        out1 => S3269
    );
nand_n_3790: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3268,
        in1(1) => S3265,
        out1 => S3271
    );
nor_n_3791: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3271,
        in1(1) => S3263,
        out1 => S3272
    );
nand_n_3792: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3269,
        in1(1) => S3262,
        out1 => S3273
    );
nor_n_3793: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3269,
        in1(1) => S3262,
        out1 => S3274
    );
nand_n_3794: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3271,
        in1(1) => S3263,
        out1 => S3275
    );
nor_n_3795: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3274,
        in1(1) => S3272,
        out1 => S3276
    );
nand_n_3796: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3275,
        in1(1) => S3273,
        out1 => S3277
    );
nor_n_3797: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3277,
        in1(1) => S3260,
        out1 => S3278
    );
nand_n_3798: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3276,
        in1(1) => S3261,
        out1 => S3279
    );
nor_n_3799: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3276,
        in1(1) => S3261,
        out1 => S3280
    );
nand_n_3800: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3277,
        in1(1) => S3260,
        out1 => S3282
    );
nor_n_3801: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3280,
        in1(1) => S3278,
        out1 => S3283
    );
nand_n_3802: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3282,
        in1(1) => S3279,
        out1 => S3284
    );
nor_n_3803: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3284,
        in1(1) => S3258,
        out1 => S3285
    );
nand_n_3804: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3283,
        in1(1) => S3257,
        out1 => S3286
    );
nor_n_3805: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3283,
        in1(1) => S3257,
        out1 => S3287
    );
nand_n_3806: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3284,
        in1(1) => S3258,
        out1 => S3288
    );
nor_n_3807: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3287,
        in1(1) => S3285,
        out1 => S3289
    );
nand_n_3808: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3288,
        in1(1) => S3286,
        out1 => S3290
    );
nor_n_3809: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3290,
        in1(1) => S3239,
        out1 => S3291
    );
nand_n_3810: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3289,
        in1(1) => S3240,
        out1 => S3293
    );
nor_n_3811: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3289,
        in1(1) => S3240,
        out1 => S3294
    );
nand_n_3812: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3290,
        in1(1) => S3239,
        out1 => S3295
    );
nor_n_3813: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3294,
        in1(1) => S3291,
        out1 => S3296
    );
nand_n_3814: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3295,
        in1(1) => S3293,
        out1 => S3297
    );
nor_n_3815: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3297,
        in1(1) => S3238,
        out1 => S3298
    );
nand_n_3816: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3296,
        in1(1) => S3236,
        out1 => S3299
    );
nor_n_3817: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3296,
        in1(1) => S3236,
        out1 => S3300
    );
nand_n_3818: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3297,
        in1(1) => S3238,
        out1 => S3301
    );
nor_n_3819: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3300,
        in1(1) => S3298,
        out1 => S3302
    );
nand_n_3820: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3301,
        in1(1) => S3299,
        out1 => S3304
    );
nor_n_3821: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3304,
        in1(1) => S3199,
        out1 => S3305
    );
nand_n_3822: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3302,
        in1(1) => S3200,
        out1 => S3306
    );
nor_n_3823: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3302,
        in1(1) => S3200,
        out1 => S3307
    );
nand_n_3824: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3304,
        in1(1) => S3199,
        out1 => S3308
    );
nor_n_3825: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3307,
        in1(1) => S3305,
        out1 => S3309
    );
nand_n_3826: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3308,
        in1(1) => S3306,
        out1 => S3310
    );
nor_n_3827: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3310,
        in1(1) => S3198,
        out1 => S3311
    );
nand_n_3828: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3309,
        in1(1) => S3197,
        out1 => S3312
    );
nor_n_3829: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3309,
        in1(1) => S3197,
        out1 => S3313
    );
nand_n_3830: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3310,
        in1(1) => S3198,
        out1 => S3315
    );
nor_n_3831: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3313,
        in1(1) => S3311,
        out1 => S3316
    );
nand_n_3832: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3315,
        in1(1) => S3312,
        out1 => S3317
    );
nor_n_3833: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3317,
        in1(1) => S3164,
        out1 => S3318
    );
nand_n_3834: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3316,
        in1(1) => S3165,
        out1 => S3319
    );
nor_n_3835: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3316,
        in1(1) => S3165,
        out1 => S3320
    );
nand_n_3836: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3317,
        in1(1) => S3164,
        out1 => S3321
    );
nor_n_3837: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3320,
        in1(1) => S3318,
        out1 => S3322
    );
nand_n_3838: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3321,
        in1(1) => S3319,
        out1 => S3323
    );
nor_n_3839: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3323,
        in1(1) => S3008,
        out1 => S3324
    );
nand_n_3840: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3322,
        in1(1) => S3006,
        out1 => S3326
    );
nand_n_3841: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3323,
        in1(1) => S3008,
        out1 => S3327
    );
nand_n_3842: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3327,
        in1(1) => S3326,
        out1 => S3328
    );
notg_3843: ENTITY WORK.notg
    PORT MAP (
        in1 => S3328,
        out1 => S3329
    );
nand_n_3844: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3328,
        in1(1) => S3162,
        out1 => S3330
    );
nand_n_3845: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3329,
        in1(1) => S3163,
        out1 => S3331
    );
notg_3846: ENTITY WORK.notg
    PORT MAP (
        in1 => S3331,
        out1 => S3332
    );
nand_n_3847: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3331,
        in1(1) => S3330,
        out1 => S3333
    );
nor_n_3848: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3333,
        in1(1) => S3142,
        out1 => S3334
    );
notg_3849: ENTITY WORK.notg
    PORT MAP (
        in1 => S3334,
        out1 => S3335
    );
nand_n_3850: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3333,
        in1(1) => S3142,
        out1 => S3337
    );
nand_n_3851: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3337,
        in1(1) => S3335,
        out1 => S3338
    );
nor_n_3852: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3338,
        in1(1) => S3161,
        out1 => S3339
    );
nand_n_3853: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3338,
        in1(1) => S3161,
        out1 => S3340
    );
nand_n_3854: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3340,
        in1(1) => S5579,
        out1 => S3341
    );
nor_n_3855: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3341,
        in1(1) => S3339,
        out1 => S3342
    );
nor_n_3856: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3342,
        in1(1) => S3158,
        out1 => S3343
    );
nand_n_3857: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3343,
        in1(1) => S3159,
        out1 => S31
    );
nor_n_3858: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3339,
        in1(1) => S3334,
        out1 => S3344
    );
nor_n_3859: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3324,
        in1(1) => S3318,
        out1 => S3345
    );
nand_n_3860: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3326,
        in1(1) => S3319,
        out1 => S3347
    );
nor_n_3861: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3311,
        in1(1) => S3305,
        out1 => S3348
    );
nand_n_3862: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3312,
        in1(1) => S3306,
        out1 => S3349
    );
nor_n_3863: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5975,
        in1(1) => S3434,
        out1 => S3350
    );
nand_n_3864: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_0,
        in1(1) => new_datapath_multdivunit_1697_B_12,
        out1 => S3351
    );
nor_n_3865: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3177,
        in1(1) => S3173,
        out1 => S3352
    );
nand_n_3866: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3178,
        in1(1) => S3174,
        out1 => S3353
    );
nand_n_3867: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_1,
        in1(1) => new_datapath_multdivunit_1697_B_11,
        out1 => S3354
    );
nand_n_3868: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_3,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S3355
    );
nand_n_3869: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3355,
        in1(1) => S3172,
        out1 => S3356
    );
nor_n_3870: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5947,
        in1(1) => S3456,
        out1 => S3358
    );
nand_n_3871: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_3,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S3359
    );
nor_n_3872: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3355,
        in1(1) => S3172,
        out1 => S3360
    );
notg_3873: ENTITY WORK.notg
    PORT MAP (
        in1 => S3360,
        out1 => S3361
    );
nand_n_3874: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3361,
        in1(1) => S3356,
        out1 => S3362
    );
nor_n_3875: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3362,
        in1(1) => S3354,
        out1 => S3363
    );
notg_3876: ENTITY WORK.notg
    PORT MAP (
        in1 => S3363,
        out1 => S3364
    );
nand_n_3877: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3362,
        in1(1) => S3354,
        out1 => S3365
    );
notg_3878: ENTITY WORK.notg
    PORT MAP (
        in1 => S3365,
        out1 => S3366
    );
nor_n_3879: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3366,
        in1(1) => S3363,
        out1 => S3367
    );
nand_n_3880: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3365,
        in1(1) => S3364,
        out1 => S3369
    );
nor_n_3881: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3369,
        in1(1) => S3352,
        out1 => S3370
    );
nand_n_3882: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3367,
        in1(1) => S3353,
        out1 => S3371
    );
nor_n_3883: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3367,
        in1(1) => S3353,
        out1 => S3372
    );
nand_n_3884: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3369,
        in1(1) => S3352,
        out1 => S3373
    );
nor_n_3885: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3372,
        in1(1) => S3370,
        out1 => S3374
    );
nand_n_3886: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3373,
        in1(1) => S3371,
        out1 => S3375
    );
nor_n_3887: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3375,
        in1(1) => S3351,
        out1 => S3376
    );
nand_n_3888: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3374,
        in1(1) => S3350,
        out1 => S3377
    );
nor_n_3889: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3374,
        in1(1) => S3350,
        out1 => S3378
    );
nand_n_3890: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3375,
        in1(1) => S3351,
        out1 => S3380
    );
nor_n_3891: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3378,
        in1(1) => S3376,
        out1 => S3381
    );
nand_n_3892: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3380,
        in1(1) => S3377,
        out1 => S3382
    );
nor_n_3893: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3234,
        in1(1) => S3225,
        out1 => S3383
    );
nand_n_3894: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3235,
        in1(1) => S3227,
        out1 => S3384
    );
nor_n_3895: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3383,
        in1(1) => S3382,
        out1 => S3385
    );
nand_n_3896: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3384,
        in1(1) => S3381,
        out1 => S3386
    );
nor_n_3897: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3384,
        in1(1) => S3381,
        out1 => S3387
    );
nand_n_3898: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3383,
        in1(1) => S3382,
        out1 => S3388
    );
nor_n_3899: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3387,
        in1(1) => S3385,
        out1 => S3389
    );
nand_n_3900: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3388,
        in1(1) => S3386,
        out1 => S3391
    );
nor_n_3901: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3391,
        in1(1) => S3185,
        out1 => S3392
    );
nand_n_3902: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3389,
        in1(1) => S3184,
        out1 => S3393
    );
nor_n_3903: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3389,
        in1(1) => S3184,
        out1 => S3394
    );
nand_n_3904: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3391,
        in1(1) => S3185,
        out1 => S3395
    );
nor_n_3905: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3394,
        in1(1) => S3392,
        out1 => S3396
    );
nand_n_3906: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3395,
        in1(1) => S3393,
        out1 => S3397
    );
nor_n_3907: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3298,
        in1(1) => S3291,
        out1 => S3398
    );
nand_n_3908: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3299,
        in1(1) => S3293,
        out1 => S3399
    );
nor_n_3909: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3217,
        in1(1) => S3212,
        out1 => S3400
    );
nand_n_3910: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3218,
        in1(1) => S3213,
        out1 => S3402
    );
nor_n_3911: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5936,
        in1(1) => S3478,
        out1 => S3403
    );
nand_n_3912: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_4,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S3404
    );
nor_n_3913: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S202,
        in1(1) => S5916,
        out1 => S3405
    );
nand_n_3914: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S203,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S3406
    );
nor_n_3915: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3405,
        in1(1) => S3210,
        out1 => S3407
    );
nand_n_3916: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3406,
        in1(1) => S3211,
        out1 => S3408
    );
nor_n_3917: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S228,
        in1(1) => S5916,
        out1 => S3409
    );
nand_n_3918: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S229,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S3410
    );
nor_n_3919: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3406,
        in1(1) => S3211,
        out1 => S3411
    );
nand_n_3920: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3405,
        in1(1) => S3210,
        out1 => S3413
    );
nor_n_3921: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3411,
        in1(1) => S3407,
        out1 => S3414
    );
nand_n_3922: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3413,
        in1(1) => S3408,
        out1 => S3415
    );
nor_n_3923: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3415,
        in1(1) => S3404,
        out1 => S3416
    );
nand_n_3924: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3414,
        in1(1) => S3403,
        out1 => S3417
    );
nor_n_3925: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3414,
        in1(1) => S3403,
        out1 => S3418
    );
nand_n_3926: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3415,
        in1(1) => S3404,
        out1 => S3419
    );
nor_n_3927: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3418,
        in1(1) => S3416,
        out1 => S3420
    );
nand_n_3928: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3419,
        in1(1) => S3417,
        out1 => S3421
    );
nor_n_3929: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3253,
        in1(1) => S3249,
        out1 => S3422
    );
nand_n_3930: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3254,
        in1(1) => S3250,
        out1 => S3424
    );
nor_n_3931: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3422,
        in1(1) => S3421,
        out1 => S3425
    );
nand_n_3932: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3424,
        in1(1) => S3420,
        out1 => S3426
    );
nor_n_3933: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3424,
        in1(1) => S3420,
        out1 => S3427
    );
nand_n_3934: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3422,
        in1(1) => S3421,
        out1 => S3428
    );
nor_n_3935: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3427,
        in1(1) => S3425,
        out1 => S3429
    );
nand_n_3936: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3428,
        in1(1) => S3426,
        out1 => S3430
    );
nor_n_3937: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3429,
        in1(1) => S3402,
        out1 => S3431
    );
nand_n_3938: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3430,
        in1(1) => S3400,
        out1 => S3432
    );
nor_n_3939: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3430,
        in1(1) => S3400,
        out1 => S3433
    );
nand_n_3940: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3429,
        in1(1) => S3402,
        out1 => S3435
    );
nor_n_3941: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3433,
        in1(1) => S3431,
        out1 => S3436
    );
nand_n_3942: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3435,
        in1(1) => S3432,
        out1 => S3437
    );
nor_n_3943: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3285,
        in1(1) => S3278,
        out1 => S3438
    );
nand_n_3944: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3286,
        in1(1) => S3279,
        out1 => S3439
    );
nor_n_3945: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S208,
        in1(1) => S5907,
        out1 => S3440
    );
nand_n_3946: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S209,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S3441
    );
nand_n_3947: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S249,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S3442
    );
nand_n_3948: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3442,
        in1(1) => S3247,
        out1 => S3443
    );
notg_3949: ENTITY WORK.notg
    PORT MAP (
        in1 => S3443,
        out1 => S3444
    );
nor_n_3950: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S240,
        in1(1) => S3336,
        out1 => S3446
    );
nand_n_3951: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S241,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S3447
    );
nor_n_3952: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3442,
        in1(1) => S3247,
        out1 => S3448
    );
nand_n_3953: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3446,
        in1(1) => S3243,
        out1 => S3449
    );
nor_n_3954: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3448,
        in1(1) => S3444,
        out1 => S3450
    );
nand_n_3955: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3449,
        in1(1) => S3443,
        out1 => S3451
    );
nor_n_3956: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3451,
        in1(1) => S3441,
        out1 => S3452
    );
nand_n_3957: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3450,
        in1(1) => S3440,
        out1 => S3453
    );
nor_n_3958: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3450,
        in1(1) => S3440,
        out1 => S3454
    );
nand_n_3959: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3451,
        in1(1) => S3441,
        out1 => S3455
    );
nor_n_3960: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3454,
        in1(1) => S3452,
        out1 => S3457
    );
nand_n_3961: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3455,
        in1(1) => S3453,
        out1 => S3458
    );
nor_n_3962: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3272,
        in1(1) => S3267,
        out1 => S3459
    );
nand_n_3963: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3273,
        in1(1) => S3268,
        out1 => S3460
    );
nand_n_3964: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S3461
    );
notg_3965: ENTITY WORK.notg
    PORT MAP (
        in1 => S3461,
        out1 => S3462
    );
nand_n_3966: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S3463
    );
nand_n_3967: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3463,
        in1(1) => S3266,
        out1 => S3464
    );
nor_n_3968: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S264,
        in1(1) => S3368,
        out1 => S3465
    );
nand_n_3969: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S265,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S3466
    );
nor_n_3970: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3466,
        in1(1) => S512,
        out1 => S3468
    );
nand_n_3971: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3465,
        in1(1) => S511,
        out1 => S3469
    );
nand_n_3972: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3469,
        in1(1) => S3464,
        out1 => S3470
    );
notg_3973: ENTITY WORK.notg
    PORT MAP (
        in1 => S3470,
        out1 => S3471
    );
nor_n_3974: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3470,
        in1(1) => S3461,
        out1 => S3472
    );
nand_n_3975: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3471,
        in1(1) => S3462,
        out1 => S3473
    );
nand_n_3976: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3470,
        in1(1) => S3461,
        out1 => S3474
    );
notg_3977: ENTITY WORK.notg
    PORT MAP (
        in1 => S3474,
        out1 => S3475
    );
nor_n_3978: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3475,
        in1(1) => S3472,
        out1 => S3476
    );
nand_n_3979: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3474,
        in1(1) => S3473,
        out1 => S3477
    );
nor_n_3980: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3477,
        in1(1) => S3459,
        out1 => S3479
    );
nand_n_3981: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3476,
        in1(1) => S3460,
        out1 => S3480
    );
nor_n_3982: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3476,
        in1(1) => S3460,
        out1 => S3481
    );
nand_n_3983: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3477,
        in1(1) => S3459,
        out1 => S3482
    );
nor_n_3984: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3481,
        in1(1) => S3479,
        out1 => S3483
    );
nand_n_3985: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3482,
        in1(1) => S3480,
        out1 => S3484
    );
nor_n_3986: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3484,
        in1(1) => S3458,
        out1 => S3485
    );
nand_n_3987: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3483,
        in1(1) => S3457,
        out1 => S3486
    );
nor_n_3988: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3483,
        in1(1) => S3457,
        out1 => S3487
    );
nand_n_3989: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3484,
        in1(1) => S3458,
        out1 => S3488
    );
nor_n_3990: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3487,
        in1(1) => S3485,
        out1 => S3490
    );
nand_n_3991: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3488,
        in1(1) => S3486,
        out1 => S3491
    );
nor_n_3992: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3491,
        in1(1) => S3438,
        out1 => S3492
    );
nand_n_3993: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3490,
        in1(1) => S3439,
        out1 => S3493
    );
nor_n_3994: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3490,
        in1(1) => S3439,
        out1 => S3494
    );
nand_n_3995: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3491,
        in1(1) => S3438,
        out1 => S3495
    );
nor_n_3996: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3494,
        in1(1) => S3492,
        out1 => S3496
    );
nand_n_3997: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3495,
        in1(1) => S3493,
        out1 => S3497
    );
nor_n_3998: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3497,
        in1(1) => S3437,
        out1 => S3498
    );
nand_n_3999: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3496,
        in1(1) => S3436,
        out1 => S3499
    );
nor_n_4000: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3496,
        in1(1) => S3436,
        out1 => S3501
    );
nand_n_4001: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3497,
        in1(1) => S3437,
        out1 => S3502
    );
nor_n_4002: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3501,
        in1(1) => S3498,
        out1 => S3503
    );
nand_n_4003: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3502,
        in1(1) => S3499,
        out1 => S3504
    );
nor_n_4004: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3504,
        in1(1) => S3398,
        out1 => S3505
    );
nand_n_4005: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3503,
        in1(1) => S3399,
        out1 => S3506
    );
nor_n_4006: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3503,
        in1(1) => S3399,
        out1 => S3507
    );
nand_n_4007: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3504,
        in1(1) => S3398,
        out1 => S3508
    );
nor_n_4008: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3507,
        in1(1) => S3505,
        out1 => S3509
    );
nand_n_4009: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3508,
        in1(1) => S3506,
        out1 => S3510
    );
nor_n_4010: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3510,
        in1(1) => S3397,
        out1 => S3512
    );
nand_n_4011: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3509,
        in1(1) => S3396,
        out1 => S3513
    );
nor_n_4012: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3509,
        in1(1) => S3396,
        out1 => S3514
    );
nand_n_4013: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3510,
        in1(1) => S3397,
        out1 => S3515
    );
nor_n_4014: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3514,
        in1(1) => S3512,
        out1 => S3516
    );
nand_n_4015: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3515,
        in1(1) => S3513,
        out1 => S3517
    );
nor_n_4016: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3517,
        in1(1) => S3348,
        out1 => S3518
    );
nand_n_4017: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3516,
        in1(1) => S3349,
        out1 => S3519
    );
nor_n_4018: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3516,
        in1(1) => S3349,
        out1 => S3520
    );
nand_n_4019: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3517,
        in1(1) => S3348,
        out1 => S3521
    );
nor_n_4020: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3520,
        in1(1) => S3518,
        out1 => S3523
    );
nand_n_4021: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3521,
        in1(1) => S3519,
        out1 => S3524
    );
nor_n_4022: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3524,
        in1(1) => S3196,
        out1 => S3525
    );
nand_n_4023: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3523,
        in1(1) => S3195,
        out1 => S3526
    );
nor_n_4024: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3523,
        in1(1) => S3195,
        out1 => S3527
    );
nand_n_4025: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3524,
        in1(1) => S3196,
        out1 => S3528
    );
nor_n_4026: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3527,
        in1(1) => S3525,
        out1 => S3529
    );
nand_n_4027: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3528,
        in1(1) => S3526,
        out1 => S3530
    );
nor_n_4028: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3529,
        in1(1) => S3347,
        out1 => S3531
    );
nand_n_4029: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3530,
        in1(1) => S3345,
        out1 => S3532
    );
nor_n_4030: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3530,
        in1(1) => S3345,
        out1 => S3534
    );
nand_n_4031: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3529,
        in1(1) => S3347,
        out1 => S3535
    );
nor_n_4032: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3534,
        in1(1) => S3531,
        out1 => S3536
    );
nand_n_4033: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3535,
        in1(1) => S3532,
        out1 => S3537
    );
nand_n_4034: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3536,
        in1(1) => S3332,
        out1 => S3538
    );
nand_n_4035: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3537,
        in1(1) => S3331,
        out1 => S3539
    );
nand_n_4036: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3539,
        in1(1) => S3538,
        out1 => S3540
    );
nor_n_4037: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3540,
        in1(1) => S3344,
        out1 => S3541
    );
notg_4038: ENTITY WORK.notg
    PORT MAP (
        in1 => S3541,
        out1 => S3542
    );
nand_n_4039: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3540,
        in1(1) => S3344,
        out1 => S3543
    );
nor_n_4040: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3541,
        in1(1) => S5590,
        out1 => S3545
    );
nand_n_4041: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3545,
        in1(1) => S3543,
        out1 => S3546
    );
nand_n_4042: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5611,
        in1(1) => new_datapath_multdivunit_outmdu1_12,
        out1 => S3547
    );
notg_4043: ENTITY WORK.notg
    PORT MAP (
        in1 => S3547,
        out1 => S3548
    );
nor_n_4044: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S393,
        in1(1) => S5547,
        out1 => S3549
    );
nor_n_4045: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3549,
        in1(1) => S3548,
        out1 => S3550
    );
nand_n_4046: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3550,
        in1(1) => S3546,
        out1 => S32
    );
nand_n_4047: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3542,
        in1(1) => S3538,
        out1 => S3551
    );
notg_4048: ENTITY WORK.notg
    PORT MAP (
        in1 => S3551,
        out1 => S3552
    );
nand_n_4049: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3526,
        in1(1) => S3519,
        out1 => S3553
    );
nor_n_4050: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3392,
        in1(1) => S3385,
        out1 => S3555
    );
nand_n_4051: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3393,
        in1(1) => S3386,
        out1 => S3556
    );
nor_n_4052: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3512,
        in1(1) => S3505,
        out1 => S3557
    );
nand_n_4053: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3513,
        in1(1) => S3506,
        out1 => S3558
    );
nor_n_4054: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3376,
        in1(1) => S3370,
        out1 => S3559
    );
nand_n_4055: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3377,
        in1(1) => S3371,
        out1 => S3560
    );
nand_n_4056: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_0,
        in1(1) => new_datapath_multdivunit_1697_B_13,
        out1 => S3561
    );
nand_n_4057: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_1,
        in1(1) => new_datapath_multdivunit_1697_B_12,
        out1 => S3562
    );
nand_n_4058: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3562,
        in1(1) => S3561,
        out1 => S3563
    );
notg_4059: ENTITY WORK.notg
    PORT MAP (
        in1 => S3563,
        out1 => S3564
    );
nand_n_4060: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_1,
        in1(1) => new_datapath_multdivunit_1697_B_13,
        out1 => S3566
    );
notg_4061: ENTITY WORK.notg
    PORT MAP (
        in1 => S3566,
        out1 => S3567
    );
nor_n_4062: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3566,
        in1(1) => S3351,
        out1 => S3568
    );
nand_n_4063: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3567,
        in1(1) => S3350,
        out1 => S3569
    );
nor_n_4064: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3568,
        in1(1) => S3564,
        out1 => S3570
    );
nand_n_4065: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3569,
        in1(1) => S3563,
        out1 => S3571
    );
nor_n_4066: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3363,
        in1(1) => S3360,
        out1 => S3572
    );
notg_4067: ENTITY WORK.notg
    PORT MAP (
        in1 => S3572,
        out1 => S3573
    );
nand_n_4068: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_2,
        in1(1) => new_datapath_multdivunit_1697_B_11,
        out1 => S3574
    );
notg_4069: ENTITY WORK.notg
    PORT MAP (
        in1 => S3574,
        out1 => S3575
    );
nor_n_4070: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5936,
        in1(1) => S3467,
        out1 => S3577
    );
nand_n_4071: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_4,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S3578
    );
nand_n_4072: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3578,
        in1(1) => S3359,
        out1 => S3579
    );
nand_n_4073: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_4,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S3580
    );
nor_n_4074: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3578,
        in1(1) => S3359,
        out1 => S3581
    );
nand_n_4075: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3577,
        in1(1) => S3358,
        out1 => S3582
    );
nand_n_4076: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3582,
        in1(1) => S3579,
        out1 => S3583
    );
notg_4077: ENTITY WORK.notg
    PORT MAP (
        in1 => S3583,
        out1 => S3584
    );
nor_n_4078: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3583,
        in1(1) => S3574,
        out1 => S3585
    );
nand_n_4079: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3584,
        in1(1) => S3575,
        out1 => S3586
    );
nand_n_4080: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3583,
        in1(1) => S3574,
        out1 => S3588
    );
nand_n_4081: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3588,
        in1(1) => S3586,
        out1 => S3589
    );
notg_4082: ENTITY WORK.notg
    PORT MAP (
        in1 => S3589,
        out1 => S3590
    );
nor_n_4083: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3589,
        in1(1) => S3572,
        out1 => S3591
    );
nand_n_4084: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3590,
        in1(1) => S3573,
        out1 => S3592
    );
nand_n_4085: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3589,
        in1(1) => S3572,
        out1 => S3593
    );
notg_4086: ENTITY WORK.notg
    PORT MAP (
        in1 => S3593,
        out1 => S3594
    );
nor_n_4087: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3594,
        in1(1) => S3591,
        out1 => S3595
    );
nand_n_4088: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3593,
        in1(1) => S3592,
        out1 => S3596
    );
nor_n_4089: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3595,
        in1(1) => S3570,
        out1 => S3597
    );
nand_n_4090: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3596,
        in1(1) => S3571,
        out1 => S3599
    );
nor_n_4091: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3596,
        in1(1) => S3571,
        out1 => S3600
    );
nand_n_4092: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3595,
        in1(1) => S3570,
        out1 => S3601
    );
nor_n_4093: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3600,
        in1(1) => S3597,
        out1 => S3602
    );
nand_n_4094: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3601,
        in1(1) => S3599,
        out1 => S3603
    );
nor_n_4095: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3433,
        in1(1) => S3425,
        out1 => S3604
    );
nand_n_4096: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3435,
        in1(1) => S3426,
        out1 => S3605
    );
nor_n_4097: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3604,
        in1(1) => S3603,
        out1 => S3606
    );
nand_n_4098: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3605,
        in1(1) => S3602,
        out1 => S3607
    );
nor_n_4099: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3605,
        in1(1) => S3602,
        out1 => S3608
    );
nand_n_4100: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3604,
        in1(1) => S3603,
        out1 => S3610
    );
nor_n_4101: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3608,
        in1(1) => S3606,
        out1 => S3611
    );
nand_n_4102: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3610,
        in1(1) => S3607,
        out1 => S3612
    );
nor_n_4103: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3611,
        in1(1) => S3560,
        out1 => S3613
    );
nand_n_4104: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3612,
        in1(1) => S3559,
        out1 => S3614
    );
nor_n_4105: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3612,
        in1(1) => S3559,
        out1 => S3615
    );
nand_n_4106: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3611,
        in1(1) => S3560,
        out1 => S3616
    );
nor_n_4107: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3615,
        in1(1) => S3613,
        out1 => S3617
    );
nand_n_4108: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3616,
        in1(1) => S3614,
        out1 => S3618
    );
nor_n_4109: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3498,
        in1(1) => S3492,
        out1 => S3619
    );
nand_n_4110: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3499,
        in1(1) => S3493,
        out1 => S3621
    );
nor_n_4111: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3416,
        in1(1) => S3411,
        out1 => S3622
    );
nand_n_4112: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3417,
        in1(1) => S3413,
        out1 => S3623
    );
nor_n_4113: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5926,
        in1(1) => S3478,
        out1 => S3624
    );
nand_n_4114: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_5,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S3625
    );
nor_n_4115: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S202,
        in1(1) => S5907,
        out1 => S3626
    );
nand_n_4116: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S203,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S3627
    );
nor_n_4117: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3626,
        in1(1) => S3409,
        out1 => S3628
    );
nand_n_4118: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3627,
        in1(1) => S3410,
        out1 => S3629
    );
nand_n_4119: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S229,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S3630
    );
nor_n_4120: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3627,
        in1(1) => S3410,
        out1 => S3632
    );
nand_n_4121: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3626,
        in1(1) => S3409,
        out1 => S3633
    );
nor_n_4122: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3632,
        in1(1) => S3628,
        out1 => S3634
    );
nand_n_4123: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3633,
        in1(1) => S3629,
        out1 => S3635
    );
nor_n_4124: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3635,
        in1(1) => S3625,
        out1 => S3636
    );
nand_n_4125: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3634,
        in1(1) => S3624,
        out1 => S3637
    );
nor_n_4126: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3634,
        in1(1) => S3624,
        out1 => S3638
    );
nand_n_4127: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3635,
        in1(1) => S3625,
        out1 => S3639
    );
nor_n_4128: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3638,
        in1(1) => S3636,
        out1 => S3640
    );
nand_n_4129: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3639,
        in1(1) => S3637,
        out1 => S3641
    );
nor_n_4130: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3452,
        in1(1) => S3448,
        out1 => S3643
    );
nand_n_4131: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3453,
        in1(1) => S3449,
        out1 => S3644
    );
nor_n_4132: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3643,
        in1(1) => S3641,
        out1 => S3645
    );
nand_n_4133: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3644,
        in1(1) => S3640,
        out1 => S3646
    );
nor_n_4134: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3644,
        in1(1) => S3640,
        out1 => S3647
    );
nand_n_4135: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3643,
        in1(1) => S3641,
        out1 => S3648
    );
nor_n_4136: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3647,
        in1(1) => S3645,
        out1 => S3649
    );
nand_n_4137: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3648,
        in1(1) => S3646,
        out1 => S3650
    );
nor_n_4138: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3649,
        in1(1) => S3623,
        out1 => S3651
    );
nand_n_4139: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3650,
        in1(1) => S3622,
        out1 => S3652
    );
nor_n_4140: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3650,
        in1(1) => S3622,
        out1 => S3654
    );
nand_n_4141: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3649,
        in1(1) => S3623,
        out1 => S3655
    );
nor_n_4142: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3654,
        in1(1) => S3651,
        out1 => S3656
    );
nand_n_4143: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3655,
        in1(1) => S3652,
        out1 => S3657
    );
nor_n_4144: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3485,
        in1(1) => S3479,
        out1 => S3658
    );
nand_n_4145: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3486,
        in1(1) => S3480,
        out1 => S3659
    );
nand_n_4146: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S209,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S3660
    );
notg_4147: ENTITY WORK.notg
    PORT MAP (
        in1 => S3660,
        out1 => S3661
    );
nor_n_4148: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S248,
        in1(1) => S3346,
        out1 => S3662
    );
nand_n_4149: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S249,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S3663
    );
nand_n_4150: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3663,
        in1(1) => S3447,
        out1 => S3665
    );
nand_n_4151: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S241,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S3666
    );
nor_n_4152: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3663,
        in1(1) => S3447,
        out1 => S3667
    );
nand_n_4153: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3662,
        in1(1) => S3446,
        out1 => S3668
    );
nand_n_4154: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3668,
        in1(1) => S3665,
        out1 => S3669
    );
notg_4155: ENTITY WORK.notg
    PORT MAP (
        in1 => S3669,
        out1 => S3670
    );
nor_n_4156: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3669,
        in1(1) => S3660,
        out1 => S3671
    );
nand_n_4157: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3670,
        in1(1) => S3661,
        out1 => S3672
    );
nand_n_4158: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3669,
        in1(1) => S3660,
        out1 => S3673
    );
notg_4159: ENTITY WORK.notg
    PORT MAP (
        in1 => S3673,
        out1 => S3674
    );
nor_n_4160: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3674,
        in1(1) => S3671,
        out1 => S3676
    );
nand_n_4161: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3673,
        in1(1) => S3672,
        out1 => S3677
    );
nor_n_4162: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3472,
        in1(1) => S3468,
        out1 => S3678
    );
nand_n_4163: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3473,
        in1(1) => S3469,
        out1 => S3679
    );
nor_n_4164: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S256,
        in1(1) => S3357,
        out1 => S3680
    );
nand_n_4165: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S3681
    );
nor_n_4166: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3465,
        in1(1) => S351,
        out1 => S3682
    );
nand_n_4167: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3466,
        in1(1) => S352,
        out1 => S3683
    );
nand_n_4168: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S265,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S3684
    );
nor_n_4169: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3466,
        in1(1) => S352,
        out1 => S3685
    );
nand_n_4170: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3465,
        in1(1) => S351,
        out1 => S3687
    );
nor_n_4171: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3685,
        in1(1) => S3682,
        out1 => S3688
    );
nand_n_4172: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3687,
        in1(1) => S3683,
        out1 => S3689
    );
nor_n_4173: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3689,
        in1(1) => S3681,
        out1 => S3690
    );
nand_n_4174: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3688,
        in1(1) => S3680,
        out1 => S3691
    );
nor_n_4175: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3688,
        in1(1) => S3680,
        out1 => S3692
    );
nand_n_4176: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3689,
        in1(1) => S3681,
        out1 => S3693
    );
nor_n_4177: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3692,
        in1(1) => S3690,
        out1 => S3694
    );
nand_n_4178: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3693,
        in1(1) => S3691,
        out1 => S3695
    );
nor_n_4179: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3695,
        in1(1) => S3678,
        out1 => S3696
    );
nand_n_4180: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3694,
        in1(1) => S3679,
        out1 => S3698
    );
nor_n_4181: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3694,
        in1(1) => S3679,
        out1 => S3699
    );
nand_n_4182: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3695,
        in1(1) => S3678,
        out1 => S3700
    );
nor_n_4183: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3699,
        in1(1) => S3696,
        out1 => S3701
    );
nand_n_4184: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3700,
        in1(1) => S3698,
        out1 => S3702
    );
nor_n_4185: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3702,
        in1(1) => S3677,
        out1 => S3703
    );
nand_n_4186: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3701,
        in1(1) => S3676,
        out1 => S3704
    );
nor_n_4187: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3701,
        in1(1) => S3676,
        out1 => S3705
    );
nand_n_4188: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3702,
        in1(1) => S3677,
        out1 => S3706
    );
nor_n_4189: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3705,
        in1(1) => S3703,
        out1 => S3707
    );
nand_n_4190: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3706,
        in1(1) => S3704,
        out1 => S3709
    );
nor_n_4191: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3709,
        in1(1) => S3658,
        out1 => S3710
    );
nand_n_4192: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3707,
        in1(1) => S3659,
        out1 => S3711
    );
nor_n_4193: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3707,
        in1(1) => S3659,
        out1 => S3712
    );
nand_n_4194: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3709,
        in1(1) => S3658,
        out1 => S3713
    );
nor_n_4195: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3712,
        in1(1) => S3710,
        out1 => S3714
    );
nand_n_4196: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3713,
        in1(1) => S3711,
        out1 => S3715
    );
nor_n_4197: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3715,
        in1(1) => S3657,
        out1 => S3716
    );
nand_n_4198: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3714,
        in1(1) => S3656,
        out1 => S3717
    );
nor_n_4199: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3714,
        in1(1) => S3656,
        out1 => S3718
    );
nand_n_4200: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3715,
        in1(1) => S3657,
        out1 => S3720
    );
nor_n_4201: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3718,
        in1(1) => S3716,
        out1 => S3721
    );
nand_n_4202: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3720,
        in1(1) => S3717,
        out1 => S3722
    );
nor_n_4203: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3722,
        in1(1) => S3619,
        out1 => S3723
    );
nand_n_4204: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3721,
        in1(1) => S3621,
        out1 => S3724
    );
nor_n_4205: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3721,
        in1(1) => S3621,
        out1 => S3725
    );
nand_n_4206: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3722,
        in1(1) => S3619,
        out1 => S3726
    );
nor_n_4207: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3725,
        in1(1) => S3723,
        out1 => S3727
    );
nand_n_4208: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3726,
        in1(1) => S3724,
        out1 => S3728
    );
nor_n_4209: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3728,
        in1(1) => S3618,
        out1 => S3729
    );
nand_n_4210: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3727,
        in1(1) => S3617,
        out1 => S3730
    );
nor_n_4211: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3727,
        in1(1) => S3617,
        out1 => S3731
    );
nand_n_4212: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3728,
        in1(1) => S3618,
        out1 => S3732
    );
nor_n_4213: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3731,
        in1(1) => S3729,
        out1 => S3733
    );
nand_n_4214: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3732,
        in1(1) => S3730,
        out1 => S3734
    );
nor_n_4215: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3734,
        in1(1) => S3557,
        out1 => S3735
    );
nand_n_4216: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3733,
        in1(1) => S3558,
        out1 => S3736
    );
nor_n_4217: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3733,
        in1(1) => S3558,
        out1 => S3737
    );
nand_n_4218: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3734,
        in1(1) => S3557,
        out1 => S3738
    );
nor_n_4219: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3737,
        in1(1) => S3735,
        out1 => S3739
    );
nand_n_4220: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3738,
        in1(1) => S3736,
        out1 => S3741
    );
nor_n_4221: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3741,
        in1(1) => S3555,
        out1 => S3742
    );
nor_n_4222: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3739,
        in1(1) => S3556,
        out1 => S3743
    );
nor_n_4223: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3743,
        in1(1) => S3742,
        out1 => S3744
    );
nor_n_4224: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3744,
        in1(1) => S3553,
        out1 => S3745
    );
notg_4225: ENTITY WORK.notg
    PORT MAP (
        in1 => S3745,
        out1 => S3746
    );
nand_n_4226: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3744,
        in1(1) => S3553,
        out1 => S3747
    );
notg_4227: ENTITY WORK.notg
    PORT MAP (
        in1 => S3747,
        out1 => S3748
    );
nor_n_4228: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3748,
        in1(1) => S3745,
        out1 => S3749
    );
nand_n_4229: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3747,
        in1(1) => S3746,
        out1 => S3750
    );
nor_n_4230: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3749,
        in1(1) => S3534,
        out1 => S3751
    );
nor_n_4231: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3750,
        in1(1) => S3535,
        out1 => S3752
    );
nor_n_4232: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3752,
        in1(1) => S3751,
        out1 => S3753
    );
nor_n_4233: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3751,
        in1(1) => S3552,
        out1 => S3754
    );
nor_n_4234: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3753,
        in1(1) => S3551,
        out1 => S3755
    );
nor_n_4235: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3755,
        in1(1) => S3754,
        out1 => S3756
    );
nand_n_4236: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3756,
        in1(1) => S5579,
        out1 => S3757
    );
nor_n_4237: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S332,
        in1(1) => S5547,
        out1 => S3758
    );
nand_n_4238: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5611,
        in1(1) => new_datapath_multdivunit_outmdu1_13,
        out1 => S3759
    );
notg_4239: ENTITY WORK.notg
    PORT MAP (
        in1 => S3759,
        out1 => S3760
    );
nor_n_4240: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3760,
        in1(1) => S3758,
        out1 => S3762
    );
nand_n_4241: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3762,
        in1(1) => S3757,
        out1 => S33
    );
nor_n_4242: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3742,
        in1(1) => S3735,
        out1 => S3763
    );
notg_4243: ENTITY WORK.notg
    PORT MAP (
        in1 => S3763,
        out1 => S3764
    );
nor_n_4244: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3615,
        in1(1) => S3606,
        out1 => S3765
    );
nand_n_4245: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3616,
        in1(1) => S3607,
        out1 => S3766
    );
nor_n_4246: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3765,
        in1(1) => S3569,
        out1 => S3767
    );
nand_n_4247: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3766,
        in1(1) => S3568,
        out1 => S3768
    );
nor_n_4248: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3766,
        in1(1) => S3568,
        out1 => S3769
    );
nand_n_4249: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3765,
        in1(1) => S3569,
        out1 => S3770
    );
nor_n_4250: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3769,
        in1(1) => S3767,
        out1 => S3772
    );
nand_n_4251: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3770,
        in1(1) => S3768,
        out1 => S3773
    );
nor_n_4252: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3729,
        in1(1) => S3723,
        out1 => S3774
    );
nand_n_4253: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3730,
        in1(1) => S3724,
        out1 => S3775
    );
nor_n_4254: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3600,
        in1(1) => S3591,
        out1 => S3776
    );
nand_n_4255: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3601,
        in1(1) => S3592,
        out1 => S3777
    );
nand_n_4256: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_0,
        in1(1) => new_datapath_multdivunit_1697_B_14,
        out1 => S3778
    );
nand_n_4257: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_2,
        in1(1) => new_datapath_multdivunit_1697_B_12,
        out1 => S3779
    );
nand_n_4258: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3779,
        in1(1) => S3566,
        out1 => S3780
    );
nor_n_4259: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5957,
        in1(1) => S3423,
        out1 => S3781
    );
nand_n_4260: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_2,
        in1(1) => new_datapath_multdivunit_1697_B_13,
        out1 => S3783
    );
nor_n_4261: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3783,
        in1(1) => S3562,
        out1 => S3784
    );
notg_4262: ENTITY WORK.notg
    PORT MAP (
        in1 => S3784,
        out1 => S3785
    );
nand_n_4263: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3785,
        in1(1) => S3780,
        out1 => S3786
    );
nor_n_4264: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3786,
        in1(1) => S3778,
        out1 => S3787
    );
notg_4265: ENTITY WORK.notg
    PORT MAP (
        in1 => S3787,
        out1 => S3788
    );
nand_n_4266: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3786,
        in1(1) => S3778,
        out1 => S3789
    );
notg_4267: ENTITY WORK.notg
    PORT MAP (
        in1 => S3789,
        out1 => S3790
    );
nor_n_4268: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3790,
        in1(1) => S3787,
        out1 => S3791
    );
nand_n_4269: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3789,
        in1(1) => S3788,
        out1 => S3792
    );
nor_n_4270: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3585,
        in1(1) => S3581,
        out1 => S3794
    );
nand_n_4271: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3586,
        in1(1) => S3582,
        out1 => S3795
    );
nand_n_4272: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_3,
        in1(1) => new_datapath_multdivunit_1697_B_11,
        out1 => S3796
    );
notg_4273: ENTITY WORK.notg
    PORT MAP (
        in1 => S3796,
        out1 => S3797
    );
nand_n_4274: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_5,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S3798
    );
nand_n_4275: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3798,
        in1(1) => S3580,
        out1 => S3799
    );
nor_n_4276: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5926,
        in1(1) => S3456,
        out1 => S3800
    );
nand_n_4277: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_5,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S3801
    );
nor_n_4278: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3801,
        in1(1) => S3578,
        out1 => S3802
    );
nand_n_4279: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3800,
        in1(1) => S3577,
        out1 => S3803
    );
nand_n_4280: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3803,
        in1(1) => S3799,
        out1 => S3805
    );
notg_4281: ENTITY WORK.notg
    PORT MAP (
        in1 => S3805,
        out1 => S3806
    );
nor_n_4282: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3805,
        in1(1) => S3796,
        out1 => S3807
    );
nand_n_4283: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3806,
        in1(1) => S3797,
        out1 => S3808
    );
nand_n_4284: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3805,
        in1(1) => S3796,
        out1 => S3809
    );
notg_4285: ENTITY WORK.notg
    PORT MAP (
        in1 => S3809,
        out1 => S3810
    );
nor_n_4286: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3810,
        in1(1) => S3807,
        out1 => S3811
    );
nand_n_4287: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3809,
        in1(1) => S3808,
        out1 => S3812
    );
nor_n_4288: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3812,
        in1(1) => S3794,
        out1 => S3813
    );
nand_n_4289: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3811,
        in1(1) => S3795,
        out1 => S3814
    );
nor_n_4290: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3811,
        in1(1) => S3795,
        out1 => S3816
    );
nand_n_4291: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3812,
        in1(1) => S3794,
        out1 => S3817
    );
nor_n_4292: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3816,
        in1(1) => S3813,
        out1 => S3818
    );
nand_n_4293: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3817,
        in1(1) => S3814,
        out1 => S3819
    );
nor_n_4294: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3818,
        in1(1) => S3791,
        out1 => S3820
    );
nand_n_4295: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3819,
        in1(1) => S3792,
        out1 => S3821
    );
nor_n_4296: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3819,
        in1(1) => S3792,
        out1 => S3822
    );
nand_n_4297: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3818,
        in1(1) => S3791,
        out1 => S3823
    );
nor_n_4298: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3822,
        in1(1) => S3820,
        out1 => S3824
    );
nand_n_4299: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3823,
        in1(1) => S3821,
        out1 => S3825
    );
nor_n_4300: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3654,
        in1(1) => S3645,
        out1 => S3827
    );
nand_n_4301: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3655,
        in1(1) => S3646,
        out1 => S3828
    );
nor_n_4302: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3827,
        in1(1) => S3825,
        out1 => S3829
    );
nand_n_4303: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3828,
        in1(1) => S3824,
        out1 => S3830
    );
nor_n_4304: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3828,
        in1(1) => S3824,
        out1 => S3831
    );
nand_n_4305: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3827,
        in1(1) => S3825,
        out1 => S3832
    );
nor_n_4306: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3831,
        in1(1) => S3829,
        out1 => S3833
    );
nand_n_4307: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3832,
        in1(1) => S3830,
        out1 => S3834
    );
nor_n_4308: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3833,
        in1(1) => S3777,
        out1 => S3835
    );
nand_n_4309: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3834,
        in1(1) => S3776,
        out1 => S3836
    );
nor_n_4310: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3834,
        in1(1) => S3776,
        out1 => S3838
    );
nand_n_4311: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3833,
        in1(1) => S3777,
        out1 => S3839
    );
nor_n_4312: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3838,
        in1(1) => S3835,
        out1 => S3840
    );
nand_n_4313: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3839,
        in1(1) => S3836,
        out1 => S3841
    );
nor_n_4314: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3716,
        in1(1) => S3710,
        out1 => S3842
    );
nand_n_4315: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3717,
        in1(1) => S3711,
        out1 => S3843
    );
nor_n_4316: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3636,
        in1(1) => S3632,
        out1 => S3844
    );
nand_n_4317: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3637,
        in1(1) => S3633,
        out1 => S3845
    );
nand_n_4318: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_6,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S3846
    );
notg_4319: ENTITY WORK.notg
    PORT MAP (
        in1 => S3846,
        out1 => S3847
    );
nand_n_4320: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S203,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S3849
    );
nand_n_4321: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3849,
        in1(1) => S3630,
        out1 => S3850
    );
nor_n_4322: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S228,
        in1(1) => S3325,
        out1 => S3851
    );
nand_n_4323: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S229,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S3852
    );
nor_n_4324: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3852,
        in1(1) => S3627,
        out1 => S3853
    );
nand_n_4325: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3851,
        in1(1) => S3626,
        out1 => S3854
    );
nand_n_4326: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3854,
        in1(1) => S3850,
        out1 => S3855
    );
notg_4327: ENTITY WORK.notg
    PORT MAP (
        in1 => S3855,
        out1 => S3856
    );
nor_n_4328: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3855,
        in1(1) => S3846,
        out1 => S3857
    );
nand_n_4329: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3856,
        in1(1) => S3847,
        out1 => S3858
    );
nand_n_4330: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3855,
        in1(1) => S3846,
        out1 => S3860
    );
notg_4331: ENTITY WORK.notg
    PORT MAP (
        in1 => S3860,
        out1 => S3861
    );
nor_n_4332: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3861,
        in1(1) => S3857,
        out1 => S3862
    );
nand_n_4333: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3860,
        in1(1) => S3858,
        out1 => S3863
    );
nor_n_4334: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3671,
        in1(1) => S3667,
        out1 => S3864
    );
nand_n_4335: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3672,
        in1(1) => S3668,
        out1 => S3865
    );
nor_n_4336: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3864,
        in1(1) => S3863,
        out1 => S3866
    );
nand_n_4337: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3865,
        in1(1) => S3862,
        out1 => S3867
    );
nor_n_4338: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3865,
        in1(1) => S3862,
        out1 => S3868
    );
nand_n_4339: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3864,
        in1(1) => S3863,
        out1 => S3869
    );
nor_n_4340: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3868,
        in1(1) => S3866,
        out1 => S3871
    );
nand_n_4341: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3869,
        in1(1) => S3867,
        out1 => S3872
    );
nor_n_4342: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3871,
        in1(1) => S3845,
        out1 => S3873
    );
nand_n_4343: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3872,
        in1(1) => S3844,
        out1 => S3874
    );
nor_n_4344: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3872,
        in1(1) => S3844,
        out1 => S3875
    );
nand_n_4345: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3871,
        in1(1) => S3845,
        out1 => S3876
    );
nor_n_4346: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3875,
        in1(1) => S3873,
        out1 => S3877
    );
nand_n_4347: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3876,
        in1(1) => S3874,
        out1 => S3878
    );
nor_n_4348: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3703,
        in1(1) => S3696,
        out1 => S3879
    );
nand_n_4349: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3704,
        in1(1) => S3698,
        out1 => S3880
    );
nand_n_4350: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S209,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S3882
    );
notg_4351: ENTITY WORK.notg
    PORT MAP (
        in1 => S3882,
        out1 => S3883
    );
nand_n_4352: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S249,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S3884
    );
nand_n_4353: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3884,
        in1(1) => S3666,
        out1 => S3885
    );
nor_n_4354: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S240,
        in1(1) => S3357,
        out1 => S3886
    );
nand_n_4355: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S241,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S3887
    );
nor_n_4356: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3887,
        in1(1) => S3663,
        out1 => S3888
    );
nand_n_4357: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3886,
        in1(1) => S3662,
        out1 => S3889
    );
nand_n_4358: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3889,
        in1(1) => S3885,
        out1 => S3890
    );
notg_4359: ENTITY WORK.notg
    PORT MAP (
        in1 => S3890,
        out1 => S3891
    );
nor_n_4360: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3890,
        in1(1) => S3882,
        out1 => S3893
    );
nand_n_4361: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3891,
        in1(1) => S3883,
        out1 => S3894
    );
nand_n_4362: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3890,
        in1(1) => S3882,
        out1 => S3895
    );
notg_4363: ENTITY WORK.notg
    PORT MAP (
        in1 => S3895,
        out1 => S3896
    );
nor_n_4364: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3896,
        in1(1) => S3893,
        out1 => S3897
    );
nand_n_4365: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3895,
        in1(1) => S3894,
        out1 => S3898
    );
nor_n_4366: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3690,
        in1(1) => S3685,
        out1 => S3899
    );
nand_n_4367: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3691,
        in1(1) => S3687,
        out1 => S3900
    );
nand_n_4368: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S3901
    );
notg_4369: ENTITY WORK.notg
    PORT MAP (
        in1 => S3901,
        out1 => S3902
    );
nand_n_4370: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S3904
    );
nand_n_4371: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3904,
        in1(1) => S3684,
        out1 => S3905
    );
nor_n_4372: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S264,
        in1(1) => S3390,
        out1 => S3906
    );
nand_n_4373: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S265,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S3907
    );
nor_n_4374: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3907,
        in1(1) => S352,
        out1 => S3908
    );
nand_n_4375: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3906,
        in1(1) => S351,
        out1 => S3909
    );
nand_n_4376: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3909,
        in1(1) => S3905,
        out1 => S3910
    );
notg_4377: ENTITY WORK.notg
    PORT MAP (
        in1 => S3910,
        out1 => S3911
    );
nor_n_4378: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3910,
        in1(1) => S3901,
        out1 => S3912
    );
nand_n_4379: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3911,
        in1(1) => S3902,
        out1 => S3913
    );
nand_n_4380: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3910,
        in1(1) => S3901,
        out1 => S3915
    );
notg_4381: ENTITY WORK.notg
    PORT MAP (
        in1 => S3915,
        out1 => S3916
    );
nor_n_4382: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3916,
        in1(1) => S3912,
        out1 => S3917
    );
nand_n_4383: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3915,
        in1(1) => S3913,
        out1 => S3918
    );
nor_n_4384: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3918,
        in1(1) => S3899,
        out1 => S3919
    );
nand_n_4385: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3917,
        in1(1) => S3900,
        out1 => S3920
    );
nor_n_4386: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3917,
        in1(1) => S3900,
        out1 => S3921
    );
nand_n_4387: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3918,
        in1(1) => S3899,
        out1 => S3922
    );
nor_n_4388: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3921,
        in1(1) => S3919,
        out1 => S3923
    );
nand_n_4389: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3922,
        in1(1) => S3920,
        out1 => S3924
    );
nor_n_4390: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3924,
        in1(1) => S3898,
        out1 => S3926
    );
nand_n_4391: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3923,
        in1(1) => S3897,
        out1 => S3927
    );
nor_n_4392: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3923,
        in1(1) => S3897,
        out1 => S3928
    );
nand_n_4393: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3924,
        in1(1) => S3898,
        out1 => S3929
    );
nor_n_4394: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3928,
        in1(1) => S3926,
        out1 => S3930
    );
nand_n_4395: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3929,
        in1(1) => S3927,
        out1 => S3931
    );
nor_n_4396: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3931,
        in1(1) => S3879,
        out1 => S3932
    );
nand_n_4397: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3930,
        in1(1) => S3880,
        out1 => S3933
    );
nor_n_4398: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3930,
        in1(1) => S3880,
        out1 => S3934
    );
nand_n_4399: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3931,
        in1(1) => S3879,
        out1 => S3935
    );
nor_n_4400: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3934,
        in1(1) => S3932,
        out1 => S3937
    );
nand_n_4401: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3935,
        in1(1) => S3933,
        out1 => S3938
    );
nor_n_4402: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3938,
        in1(1) => S3878,
        out1 => S3939
    );
nand_n_4403: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3937,
        in1(1) => S3877,
        out1 => S3940
    );
nor_n_4404: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3937,
        in1(1) => S3877,
        out1 => S3941
    );
nand_n_4405: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3938,
        in1(1) => S3878,
        out1 => S3942
    );
nor_n_4406: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3941,
        in1(1) => S3939,
        out1 => S3943
    );
nand_n_4407: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3942,
        in1(1) => S3940,
        out1 => S3944
    );
nor_n_4408: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3944,
        in1(1) => S3842,
        out1 => S3945
    );
nand_n_4409: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3943,
        in1(1) => S3843,
        out1 => S3946
    );
nor_n_4410: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3943,
        in1(1) => S3843,
        out1 => S3948
    );
nand_n_4411: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3944,
        in1(1) => S3842,
        out1 => S3949
    );
nor_n_4412: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3948,
        in1(1) => S3945,
        out1 => S3950
    );
nand_n_4413: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3949,
        in1(1) => S3946,
        out1 => S3951
    );
nor_n_4414: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3951,
        in1(1) => S3841,
        out1 => S3952
    );
nand_n_4415: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3950,
        in1(1) => S3840,
        out1 => S3953
    );
nor_n_4416: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3950,
        in1(1) => S3840,
        out1 => S3954
    );
nand_n_4417: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3951,
        in1(1) => S3841,
        out1 => S3955
    );
nor_n_4418: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3954,
        in1(1) => S3952,
        out1 => S3956
    );
nand_n_4419: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3955,
        in1(1) => S3953,
        out1 => S3957
    );
nor_n_4420: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3957,
        in1(1) => S3774,
        out1 => S3959
    );
nand_n_4421: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3956,
        in1(1) => S3775,
        out1 => S3960
    );
nor_n_4422: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3956,
        in1(1) => S3775,
        out1 => S3961
    );
nand_n_4423: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3957,
        in1(1) => S3774,
        out1 => S3962
    );
nor_n_4424: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3961,
        in1(1) => S3959,
        out1 => S3963
    );
nand_n_4425: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3962,
        in1(1) => S3960,
        out1 => S3964
    );
nor_n_4426: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3964,
        in1(1) => S3773,
        out1 => S3965
    );
nand_n_4427: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3963,
        in1(1) => S3772,
        out1 => S3966
    );
nand_n_4428: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3964,
        in1(1) => S3773,
        out1 => S3967
    );
nand_n_4429: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3967,
        in1(1) => S3966,
        out1 => S3968
    );
notg_4430: ENTITY WORK.notg
    PORT MAP (
        in1 => S3968,
        out1 => S3970
    );
nand_n_4431: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3968,
        in1(1) => S3763,
        out1 => S3971
    );
nand_n_4432: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3970,
        in1(1) => S3764,
        out1 => S3972
    );
nand_n_4433: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3972,
        in1(1) => S3971,
        out1 => S3973
    );
nor_n_4434: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3973,
        in1(1) => S3747,
        out1 => S3974
    );
notg_4435: ENTITY WORK.notg
    PORT MAP (
        in1 => S3974,
        out1 => S3975
    );
nand_n_4436: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3973,
        in1(1) => S3747,
        out1 => S3976
    );
nand_n_4437: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3976,
        in1(1) => S3975,
        out1 => S3977
    );
nor_n_4438: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3754,
        in1(1) => S3752,
        out1 => S3978
    );
nor_n_4439: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3978,
        in1(1) => S3977,
        out1 => S3979
    );
nand_n_4440: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3978,
        in1(1) => S3977,
        out1 => S3981
    );
nor_n_4441: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3979,
        in1(1) => S5590,
        out1 => S3982
    );
nand_n_4442: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3982,
        in1(1) => S3981,
        out1 => S3983
    );
nand_n_4443: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5611,
        in1(1) => new_datapath_multdivunit_outmdu1_14,
        out1 => S3984
    );
notg_4444: ENTITY WORK.notg
    PORT MAP (
        in1 => S3984,
        out1 => S3985
    );
nor_n_4445: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S291,
        in1(1) => S5547,
        out1 => S3986
    );
nor_n_4446: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3986,
        in1(1) => S3985,
        out1 => S3987
    );
nand_n_4447: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3987,
        in1(1) => S3983,
        out1 => S34
    );
nor_n_4448: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3979,
        in1(1) => S3974,
        out1 => S3988
    );
nor_n_4449: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3965,
        in1(1) => S3959,
        out1 => S3989
    );
nand_n_4450: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3966,
        in1(1) => S3960,
        out1 => S3991
    );
nor_n_4451: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3822,
        in1(1) => S3813,
        out1 => S3992
    );
nand_n_4452: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3823,
        in1(1) => S3814,
        out1 => S3993
    );
nor_n_4453: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3939,
        in1(1) => S3932,
        out1 => S3994
    );
nand_n_4454: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3940,
        in1(1) => S3933,
        out1 => S3995
    );
nor_n_4455: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3995,
        in1(1) => S3992,
        out1 => S3996
    );
nand_n_4456: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3994,
        in1(1) => S3993,
        out1 => S3997
    );
nor_n_4457: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3994,
        in1(1) => S3993,
        out1 => S3998
    );
nand_n_4458: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3995,
        in1(1) => S3992,
        out1 => S3999
    );
nor_n_4459: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3998,
        in1(1) => S3996,
        out1 => S4000
    );
nand_n_4460: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3999,
        in1(1) => S3997,
        out1 => S4002
    );
nor_n_4461: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3952,
        in1(1) => S3945,
        out1 => S4003
    );
nand_n_4462: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3953,
        in1(1) => S3946,
        out1 => S4004
    );
nor_n_4463: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3875,
        in1(1) => S3866,
        out1 => S4005
    );
nand_n_4464: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3876,
        in1(1) => S3867,
        out1 => S4006
    );
nor_n_4465: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3807,
        in1(1) => S3802,
        out1 => S4007
    );
nand_n_4466: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3808,
        in1(1) => S3803,
        out1 => S4008
    );
nor_n_4467: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5936,
        in1(1) => S3445,
        out1 => S4009
    );
nand_n_4468: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_4,
        in1(1) => new_datapath_multdivunit_1697_B_11,
        out1 => S4010
    );
nor_n_4469: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5916,
        in1(1) => S3467,
        out1 => S4011
    );
nand_n_4470: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_6,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S4013
    );
nor_n_4471: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4013,
        in1(1) => S3800,
        out1 => S4014
    );
nand_n_4472: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4011,
        in1(1) => S3801,
        out1 => S4015
    );
nor_n_4473: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4011,
        in1(1) => S3801,
        out1 => S4016
    );
nand_n_4474: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4013,
        in1(1) => S3800,
        out1 => S4017
    );
nor_n_4475: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4016,
        in1(1) => S4014,
        out1 => S4018
    );
nand_n_4476: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4017,
        in1(1) => S4015,
        out1 => S4019
    );
nor_n_4477: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4019,
        in1(1) => S4010,
        out1 => S4020
    );
nand_n_4478: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4018,
        in1(1) => S4009,
        out1 => S4021
    );
nor_n_4479: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4018,
        in1(1) => S4009,
        out1 => S4022
    );
nand_n_4480: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4019,
        in1(1) => S4010,
        out1 => S4024
    );
nor_n_4481: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4022,
        in1(1) => S4020,
        out1 => S4025
    );
nand_n_4482: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4024,
        in1(1) => S4021,
        out1 => S4026
    );
nor_n_4483: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4026,
        in1(1) => S4007,
        out1 => S4027
    );
nand_n_4484: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4025,
        in1(1) => S4008,
        out1 => S4028
    );
nor_n_4485: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4025,
        in1(1) => S4008,
        out1 => S4029
    );
nand_n_4486: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4026,
        in1(1) => S4007,
        out1 => S4030
    );
nor_n_4487: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4029,
        in1(1) => S4027,
        out1 => S4031
    );
nand_n_4488: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4030,
        in1(1) => S4028,
        out1 => S4032
    );
nor_n_4489: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4032,
        in1(1) => S4006,
        out1 => S4033
    );
nand_n_4490: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4031,
        in1(1) => S4005,
        out1 => S4035
    );
nor_n_4491: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4031,
        in1(1) => S4005,
        out1 => S4036
    );
nand_n_4492: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4032,
        in1(1) => S4006,
        out1 => S4037
    );
nor_n_4493: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4036,
        in1(1) => S4033,
        out1 => S4038
    );
nand_n_4494: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4037,
        in1(1) => S4035,
        out1 => S4039
    );
nor_n_4495: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S248,
        in1(1) => S3368,
        out1 => S4040
    );
nand_n_4496: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S249,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S4041
    );
nor_n_4497: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => S3401,
        out1 => S4042
    );
nand_n_4498: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S4043
    );
nor_n_4499: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4043,
        in1(1) => S3906,
        out1 => S4044
    );
nand_n_4500: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4042,
        in1(1) => S3907,
        out1 => S4046
    );
nor_n_4501: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4042,
        in1(1) => S3907,
        out1 => S4047
    );
nand_n_4502: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4043,
        in1(1) => S3906,
        out1 => S4048
    );
nor_n_4503: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4047,
        in1(1) => S4044,
        out1 => S4049
    );
nand_n_4504: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4048,
        in1(1) => S4046,
        out1 => S4050
    );
nor_n_4505: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S208,
        in1(1) => S3346,
        out1 => S4051
    );
nand_n_4506: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S209,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S4052
    );
nor_n_4507: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S256,
        in1(1) => S3379,
        out1 => S4053
    );
nand_n_4508: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S4054
    );
nor_n_4509: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3912,
        in1(1) => S3908,
        out1 => S4055
    );
nand_n_4510: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3913,
        in1(1) => S3909,
        out1 => S4057
    );
nor_n_4511: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4041,
        in1(1) => S3886,
        out1 => S4058
    );
nand_n_4512: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4040,
        in1(1) => S3887,
        out1 => S4059
    );
nor_n_4513: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4040,
        in1(1) => S3887,
        out1 => S4060
    );
nand_n_4514: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4041,
        in1(1) => S3886,
        out1 => S4061
    );
nor_n_4515: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4060,
        in1(1) => S4058,
        out1 => S4062
    );
nand_n_4516: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4061,
        in1(1) => S4059,
        out1 => S4063
    );
nor_n_4517: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4063,
        in1(1) => S4052,
        out1 => S4064
    );
nand_n_4518: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4062,
        in1(1) => S4051,
        out1 => S4065
    );
nor_n_4519: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4062,
        in1(1) => S4051,
        out1 => S4066
    );
nand_n_4520: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4063,
        in1(1) => S4052,
        out1 => S4068
    );
nor_n_4521: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4066,
        in1(1) => S4064,
        out1 => S4069
    );
nand_n_4522: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4068,
        in1(1) => S4065,
        out1 => S4070
    );
nor_n_4523: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4054,
        in1(1) => S4050,
        out1 => S4071
    );
nand_n_4524: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4053,
        in1(1) => S4049,
        out1 => S4072
    );
nor_n_4525: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4053,
        in1(1) => S4049,
        out1 => S4073
    );
nand_n_4526: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4054,
        in1(1) => S4050,
        out1 => S4074
    );
nor_n_4527: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4073,
        in1(1) => S4071,
        out1 => S4075
    );
nand_n_4528: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4074,
        in1(1) => S4072,
        out1 => S4076
    );
nor_n_4529: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4075,
        in1(1) => S4055,
        out1 => S4077
    );
nand_n_4530: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4076,
        in1(1) => S4057,
        out1 => S4079
    );
nor_n_4531: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4076,
        in1(1) => S4057,
        out1 => S4080
    );
nand_n_4532: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4075,
        in1(1) => S4055,
        out1 => S4081
    );
nor_n_4533: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4080,
        in1(1) => S4077,
        out1 => S4082
    );
nand_n_4534: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4081,
        in1(1) => S4079,
        out1 => S4083
    );
nor_n_4535: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4083,
        in1(1) => S4069,
        out1 => S4084
    );
nand_n_4536: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4082,
        in1(1) => S4070,
        out1 => S4085
    );
nor_n_4537: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4082,
        in1(1) => S4070,
        out1 => S4086
    );
nand_n_4538: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4083,
        in1(1) => S4069,
        out1 => S4087
    );
nor_n_4539: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4086,
        in1(1) => S4084,
        out1 => S4088
    );
nand_n_4540: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4087,
        in1(1) => S4085,
        out1 => S4090
    );
nor_n_4541: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5907,
        in1(1) => S3478,
        out1 => S4091
    );
nand_n_4542: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_7,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S4092
    );
nor_n_4543: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3893,
        in1(1) => S3888,
        out1 => S4093
    );
nand_n_4544: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3894,
        in1(1) => S3889,
        out1 => S4094
    );
nor_n_4545: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S202,
        in1(1) => S3336,
        out1 => S4095
    );
nand_n_4546: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S203,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S4096
    );
nor_n_4547: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4096,
        in1(1) => S3851,
        out1 => S4097
    );
nand_n_4548: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4095,
        in1(1) => S3852,
        out1 => S4098
    );
nor_n_4549: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4095,
        in1(1) => S3852,
        out1 => S4099
    );
nand_n_4550: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4096,
        in1(1) => S3851,
        out1 => S4101
    );
nor_n_4551: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4099,
        in1(1) => S4097,
        out1 => S4102
    );
nand_n_4552: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4101,
        in1(1) => S4098,
        out1 => S4103
    );
nor_n_4553: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4103,
        in1(1) => S4094,
        out1 => S4104
    );
nand_n_4554: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4102,
        in1(1) => S4093,
        out1 => S4105
    );
nor_n_4555: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4102,
        in1(1) => S4093,
        out1 => S4106
    );
nand_n_4556: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4103,
        in1(1) => S4094,
        out1 => S4107
    );
nor_n_4557: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4106,
        in1(1) => S4104,
        out1 => S4108
    );
nand_n_4558: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4107,
        in1(1) => S4105,
        out1 => S4109
    );
nor_n_4559: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4109,
        in1(1) => S4091,
        out1 => S4110
    );
nand_n_4560: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4108,
        in1(1) => S4092,
        out1 => S4112
    );
nor_n_4561: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4108,
        in1(1) => S4092,
        out1 => S4113
    );
nand_n_4562: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4109,
        in1(1) => S4091,
        out1 => S4114
    );
nor_n_4563: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4113,
        in1(1) => S4110,
        out1 => S4115
    );
nand_n_4564: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4114,
        in1(1) => S4112,
        out1 => S4116
    );
nor_n_4565: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4116,
        in1(1) => S4090,
        out1 => S4117
    );
nand_n_4566: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4115,
        in1(1) => S4088,
        out1 => S4118
    );
nor_n_4567: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4115,
        in1(1) => S4088,
        out1 => S4119
    );
nand_n_4568: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4116,
        in1(1) => S4090,
        out1 => S4120
    );
nor_n_4569: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4119,
        in1(1) => S4117,
        out1 => S4121
    );
nand_n_4570: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4120,
        in1(1) => S4118,
        out1 => S4123
    );
nand_n_4571: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_0,
        in1(1) => new_datapath_multdivunit_1697_B_15,
        out1 => S4124
    );
nor_n_4572: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5966,
        in1(1) => S3412,
        out1 => S4125
    );
nand_n_4573: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_1,
        in1(1) => new_datapath_multdivunit_1697_B_14,
        out1 => S4126
    );
nor_n_4574: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5947,
        in1(1) => S3434,
        out1 => S4127
    );
nand_n_4575: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_3,
        in1(1) => new_datapath_multdivunit_1697_B_12,
        out1 => S4128
    );
nor_n_4576: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4128,
        in1(1) => S3781,
        out1 => S4129
    );
nand_n_4577: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4127,
        in1(1) => S3783,
        out1 => S4130
    );
nor_n_4578: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4127,
        in1(1) => S3783,
        out1 => S4131
    );
nand_n_4579: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4128,
        in1(1) => S3781,
        out1 => S4132
    );
nor_n_4580: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4131,
        in1(1) => S4129,
        out1 => S4134
    );
nand_n_4581: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4132,
        in1(1) => S4130,
        out1 => S4135
    );
nor_n_4582: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4135,
        in1(1) => S4126,
        out1 => S4136
    );
nand_n_4583: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4134,
        in1(1) => S4125,
        out1 => S4137
    );
nor_n_4584: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4134,
        in1(1) => S4125,
        out1 => S4138
    );
nand_n_4585: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4135,
        in1(1) => S4126,
        out1 => S4139
    );
nor_n_4586: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4138,
        in1(1) => S4136,
        out1 => S4140
    );
nand_n_4587: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4139,
        in1(1) => S4137,
        out1 => S4141
    );
nor_n_4588: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3787,
        in1(1) => S3784,
        out1 => S4142
    );
nor_n_4589: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3857,
        in1(1) => S3853,
        out1 => S4143
    );
nand_n_4590: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3858,
        in1(1) => S3854,
        out1 => S4145
    );
nor_n_4591: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3926,
        in1(1) => S3919,
        out1 => S4146
    );
nand_n_4592: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3927,
        in1(1) => S3920,
        out1 => S4147
    );
nor_n_4593: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4147,
        in1(1) => S4143,
        out1 => S4148
    );
nand_n_4594: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4146,
        in1(1) => S4145,
        out1 => S4149
    );
nor_n_4595: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4146,
        in1(1) => S4145,
        out1 => S4150
    );
nand_n_4596: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4147,
        in1(1) => S4143,
        out1 => S4151
    );
nor_n_4597: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4150,
        in1(1) => S4148,
        out1 => S4152
    );
nand_n_4598: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4151,
        in1(1) => S4149,
        out1 => S4153
    );
nor_n_4599: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4153,
        in1(1) => S4123,
        out1 => S4154
    );
nand_n_4600: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4152,
        in1(1) => S4121,
        out1 => S4156
    );
nor_n_4601: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4152,
        in1(1) => S4121,
        out1 => S4157
    );
nand_n_4602: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4153,
        in1(1) => S4123,
        out1 => S4158
    );
nor_n_4603: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4157,
        in1(1) => S4154,
        out1 => S4159
    );
nand_n_4604: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4158,
        in1(1) => S4156,
        out1 => S4160
    );
nand_n_4605: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4142,
        in1(1) => S4124,
        out1 => S4161
    );
notg_4606: ENTITY WORK.notg
    PORT MAP (
        in1 => S4161,
        out1 => S4162
    );
nor_n_4607: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4142,
        in1(1) => S4124,
        out1 => S4163
    );
notg_4608: ENTITY WORK.notg
    PORT MAP (
        in1 => S4163,
        out1 => S4164
    );
nor_n_4609: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4163,
        in1(1) => S4162,
        out1 => S4165
    );
nand_n_4610: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4164,
        in1(1) => S4161,
        out1 => S4167
    );
nor_n_4611: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4167,
        in1(1) => S4140,
        out1 => S4168
    );
nand_n_4612: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4165,
        in1(1) => S4141,
        out1 => S4169
    );
nor_n_4613: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4165,
        in1(1) => S4141,
        out1 => S4170
    );
nand_n_4614: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4167,
        in1(1) => S4140,
        out1 => S4171
    );
nor_n_4615: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4170,
        in1(1) => S4168,
        out1 => S4172
    );
nand_n_4616: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4171,
        in1(1) => S4169,
        out1 => S4173
    );
nor_n_4617: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4172,
        in1(1) => S4160,
        out1 => S4174
    );
nand_n_4618: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4173,
        in1(1) => S4159,
        out1 => S4175
    );
nor_n_4619: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4173,
        in1(1) => S4159,
        out1 => S4176
    );
nand_n_4620: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4172,
        in1(1) => S4160,
        out1 => S4178
    );
nor_n_4621: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4176,
        in1(1) => S4174,
        out1 => S4179
    );
nand_n_4622: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4178,
        in1(1) => S4175,
        out1 => S4180
    );
nor_n_4623: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4180,
        in1(1) => S4039,
        out1 => S4181
    );
nand_n_4624: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4179,
        in1(1) => S4038,
        out1 => S4182
    );
nor_n_4625: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4179,
        in1(1) => S4038,
        out1 => S4183
    );
nand_n_4626: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4180,
        in1(1) => S4039,
        out1 => S4184
    );
nor_n_4627: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4183,
        in1(1) => S4181,
        out1 => S4185
    );
nand_n_4628: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4184,
        in1(1) => S4182,
        out1 => S4186
    );
nor_n_4629: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3838,
        in1(1) => S3829,
        out1 => S4187
    );
nand_n_4630: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3839,
        in1(1) => S3830,
        out1 => S4189
    );
nor_n_4631: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4187,
        in1(1) => S4186,
        out1 => S4190
    );
nand_n_4632: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4189,
        in1(1) => S4185,
        out1 => S4191
    );
nor_n_4633: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4189,
        in1(1) => S4185,
        out1 => S4192
    );
nand_n_4634: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4187,
        in1(1) => S4186,
        out1 => S4193
    );
nor_n_4635: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4192,
        in1(1) => S4190,
        out1 => S4194
    );
nand_n_4636: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4193,
        in1(1) => S4191,
        out1 => S4195
    );
nor_n_4637: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4194,
        in1(1) => S4004,
        out1 => S4196
    );
nand_n_4638: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4195,
        in1(1) => S4003,
        out1 => S4197
    );
nor_n_4639: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4195,
        in1(1) => S4003,
        out1 => S4198
    );
nand_n_4640: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4194,
        in1(1) => S4004,
        out1 => S4200
    );
nor_n_4641: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4198,
        in1(1) => S4196,
        out1 => S4201
    );
nand_n_4642: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4200,
        in1(1) => S4197,
        out1 => S4202
    );
nor_n_4643: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4201,
        in1(1) => S4000,
        out1 => S4203
    );
nand_n_4644: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4202,
        in1(1) => S4002,
        out1 => S4204
    );
nor_n_4645: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4202,
        in1(1) => S4002,
        out1 => S4205
    );
nand_n_4646: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4201,
        in1(1) => S4000,
        out1 => S4206
    );
nor_n_4647: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4205,
        in1(1) => S4203,
        out1 => S4207
    );
nand_n_4648: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4206,
        in1(1) => S4204,
        out1 => S4208
    );
nor_n_4649: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4208,
        in1(1) => S3989,
        out1 => S4209
    );
nand_n_4650: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4207,
        in1(1) => S3991,
        out1 => S4211
    );
nor_n_4651: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4207,
        in1(1) => S3991,
        out1 => S4212
    );
nand_n_4652: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4208,
        in1(1) => S3989,
        out1 => S4213
    );
nor_n_4653: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4212,
        in1(1) => S4209,
        out1 => S4214
    );
nand_n_4654: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4213,
        in1(1) => S4211,
        out1 => S4215
    );
nor_n_4655: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3972,
        in1(1) => S3768,
        out1 => S4216
    );
notg_4656: ENTITY WORK.notg
    PORT MAP (
        in1 => S4216,
        out1 => S4217
    );
nand_n_4657: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3972,
        in1(1) => S3768,
        out1 => S4218
    );
notg_4658: ENTITY WORK.notg
    PORT MAP (
        in1 => S4218,
        out1 => S4219
    );
nand_n_4659: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4218,
        in1(1) => S4217,
        out1 => S4220
    );
nor_n_4660: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4219,
        in1(1) => S4216,
        out1 => S4222
    );
nand_n_4661: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4222,
        in1(1) => S4214,
        out1 => S4223
    );
nand_n_4662: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4220,
        in1(1) => S4215,
        out1 => S4224
    );
nand_n_4663: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4224,
        in1(1) => S4223,
        out1 => S4225
    );
nor_n_4664: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4225,
        in1(1) => S3988,
        out1 => S4226
    );
nand_n_4665: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4225,
        in1(1) => S3988,
        out1 => S4227
    );
nand_n_4666: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4227,
        in1(1) => S5579,
        out1 => S4228
    );
nor_n_4667: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4228,
        in1(1) => S4226,
        out1 => S4229
    );
nand_n_4668: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5611,
        in1(1) => new_datapath_multdivunit_outmdu1_15,
        out1 => S4230
    );
nor_n_4669: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S4231
    );
nor_n_4670: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4231,
        in1(1) => S5547,
        out1 => S4233
    );
nand_n_4671: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4233,
        in1(1) => S272,
        out1 => S4234
    );
nand_n_4672: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4234,
        in1(1) => S4230,
        out1 => S4235
    );
nor_n_4673: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4235,
        in1(1) => S4229,
        out1 => S4236
    );
notg_4674: ENTITY WORK.notg
    PORT MAP (
        in1 => S4236,
        out1 => S35
    );
nor_n_4675: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => S2800,
        out1 => S36
    );
nor_n_4676: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => S2811,
        out1 => S37
    );
nor_n_4677: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => S2822,
        out1 => S38
    );
nor_n_4678: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => S2832,
        out1 => S39
    );
nor_n_4679: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => S2843,
        out1 => S40
    );
nor_n_4680: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => S2854,
        out1 => S41
    );
nor_n_4681: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => S2865,
        out1 => S42
    );
nor_n_4682: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => S2876,
        out1 => S43
    );
nor_n_4683: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => S2887,
        out1 => S44
    );
nor_n_4684: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => S2898,
        out1 => S45
    );
nor_n_4685: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => S2909,
        out1 => S46
    );
nor_n_4686: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => S2920,
        out1 => S47
    );
nor_n_4687: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => S2931,
        out1 => S48
    );
nor_n_4688: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => S2942,
        out1 => S49
    );
nor_n_4689: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => S2953,
        out1 => S50
    );
nand_n_4690: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_databusin_0,
        out1 => S4239
    );
nand_n_4691: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6087,
        in1(1) => new_datapath_instruction_0,
        out1 => S4240
    );
nand_n_4692: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4240,
        in1(1) => S4239,
        out1 => S51
    );
nand_n_4693: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_databusin_1,
        out1 => S4241
    );
nand_n_4694: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6087,
        in1(1) => new_datapath_instruction_1,
        out1 => S4242
    );
nand_n_4695: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4242,
        in1(1) => S4241,
        out1 => S52
    );
nand_n_4696: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_databusin_2,
        out1 => S4243
    );
nand_n_4697: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6087,
        in1(1) => new_datapath_instruction_2,
        out1 => S4244
    );
nand_n_4698: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4244,
        in1(1) => S4243,
        out1 => S53
    );
nand_n_4699: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_databusin_3,
        out1 => S4245
    );
nand_n_4700: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6087,
        in1(1) => new_datapath_instruction_3,
        out1 => S4247
    );
nand_n_4701: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4247,
        in1(1) => S4245,
        out1 => S54
    );
nand_n_4702: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_databusin_4,
        out1 => S4248
    );
nand_n_4703: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6087,
        in1(1) => new_controller_fib_0,
        out1 => S4249
    );
nand_n_4704: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4249,
        in1(1) => S4248,
        out1 => S55
    );
nand_n_4705: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_databusin_5,
        out1 => S4250
    );
nand_n_4706: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6087,
        in1(1) => new_controller_fib_1,
        out1 => S4251
    );
nand_n_4707: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4251,
        in1(1) => S4250,
        out1 => S56
    );
nand_n_4708: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_databusin_6,
        out1 => S4252
    );
nand_n_4709: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6087,
        in1(1) => new_controller_fib_2,
        out1 => S4253
    );
nand_n_4710: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4253,
        in1(1) => S4252,
        out1 => S57
    );
nand_n_4711: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_databusin_7,
        out1 => S4255
    );
nand_n_4712: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6087,
        in1(1) => new_controller_fib_3,
        out1 => S4256
    );
nand_n_4713: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4256,
        in1(1) => S4255,
        out1 => S58
    );
nand_n_4714: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_databusin_8,
        out1 => S4257
    );
nand_n_4715: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6087,
        in1(1) => new_controller_fib_4,
        out1 => S4258
    );
nand_n_4716: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4258,
        in1(1) => S4257,
        out1 => S59
    );
nand_n_4717: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_databusin_9,
        out1 => S4259
    );
nand_n_4718: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6087,
        in1(1) => new_controller_234_B_0,
        out1 => S4260
    );
nand_n_4719: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4260,
        in1(1) => S4259,
        out1 => S60
    );
nand_n_4720: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_databusin_10,
        out1 => S4262
    );
nand_n_4721: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6087,
        in1(1) => new_controller_opcode_2,
        out1 => S4263
    );
nand_n_4722: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4263,
        in1(1) => S4262,
        out1 => S61
    );
nand_n_4723: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_databusin_11,
        out1 => S4264
    );
nand_n_4724: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6087,
        in1(1) => new_controller_opcode_3,
        out1 => S4265
    );
nand_n_4725: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4265,
        in1(1) => S4264,
        out1 => S62
    );
nand_n_4726: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_databusin_12,
        out1 => S4266
    );
nand_n_4727: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6087,
        in1(1) => new_controller_opcode_4,
        out1 => S4267
    );
nand_n_4728: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4267,
        in1(1) => S4266,
        out1 => S63
    );
nand_n_4729: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_databusin_13,
        out1 => S4268
    );
nand_n_4730: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6087,
        in1(1) => new_controller_opcode_5,
        out1 => S4270
    );
nand_n_4731: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4270,
        in1(1) => S4268,
        out1 => S64
    );
nand_n_4732: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_databusin_14,
        out1 => S4271
    );
nand_n_4733: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6087,
        in1(1) => new_controller_opcode_6,
        out1 => S4272
    );
nand_n_4734: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4272,
        in1(1) => S4271,
        out1 => S65
    );
nor_n_4735: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S172,
        in1(1) => new_controller_opcode_2,
        out1 => S4273
    );
nand_n_4736: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S171,
        in1(1) => S3051,
        out1 => S4274
    );
nand_n_4737: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4274,
        in1(1) => new_controller_407_B_0,
        out1 => S4275
    );
nor_n_4738: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4274,
        in1(1) => S3040,
        out1 => S4276
    );
nand_n_4739: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4273,
        in1(1) => new_controller_234_B_0,
        out1 => S4277
    );
nor_n_4740: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4276,
        in1(1) => S5365,
        out1 => S4279
    );
nand_n_4741: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4277,
        in1(1) => S5354,
        out1 => S4280
    );
nand_n_4742: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_2,
        in1(1) => S5157,
        out1 => S4281
    );
nor_n_4743: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5147,
        in1(1) => S4067,
        out1 => S4282
    );
nand_n_4744: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4282,
        in1(1) => S3761,
        out1 => S4283
    );
notg_4745: ENTITY WORK.notg
    PORT MAP (
        in1 => S4283,
        out1 => S4284
    );
nand_n_4746: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4283,
        in1(1) => S5343,
        out1 => S4285
    );
nand_n_4747: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4283,
        in1(1) => S5354,
        out1 => S4286
    );
nor_n_4748: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4284,
        in1(1) => S4289,
        out1 => S4287
    );
nand_n_4749: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4287,
        in1(1) => S4279,
        out1 => S4288
    );
nand_n_4750: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4288,
        in1(1) => new_controller_fib_2,
        out1 => S4290
    );
nand_n_4751: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4290,
        in1(1) => S4281,
        out1 => S4291
    );
nand_n_4752: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4291,
        in1(1) => S4280,
        out1 => S4292
    );
nor_n_4753: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S175,
        in1(1) => S5515,
        out1 => S4293
    );
nand_n_4754: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S176,
        in1(1) => S5526,
        out1 => S4294
    );
nand_n_4755: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4294,
        in1(1) => S257,
        out1 => S4295
    );
nand_n_4756: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4295,
        in1(1) => S4292,
        out1 => S4296
    );
nor_n_4757: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4296,
        in1(1) => S5957,
        out1 => S4297
    );
nand_n_4758: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4296,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S4298
    );
notg_4759: ENTITY WORK.notg
    PORT MAP (
        in1 => S4298,
        out1 => S4299
    );
nor_n_4760: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4296,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S4301
    );
nor_n_4761: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4301,
        in1(1) => S4299,
        out1 => S4302
    );
nor_n_4762: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5907,
        in1(1) => S5168,
        out1 => S4303
    );
nand_n_4763: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4286,
        in1(1) => new_controller_opcode_3,
        out1 => S4304
    );
nand_n_4764: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4276,
        in1(1) => new_controller_fib_4,
        out1 => S4305
    );
nand_n_4765: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4305,
        in1(1) => S4300,
        out1 => S4306
    );
notg_4766: ENTITY WORK.notg
    PORT MAP (
        in1 => S4306,
        out1 => S4307
    );
nor_n_4767: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4306,
        in1(1) => S4303,
        out1 => S4308
    );
nand_n_4768: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4308,
        in1(1) => S4304,
        out1 => S4309
    );
nand_n_4769: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4309,
        in1(1) => S4280,
        out1 => S4310
    );
nand_n_4770: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4294,
        in1(1) => S229,
        out1 => S4312
    );
nand_n_4771: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4312,
        in1(1) => S4310,
        out1 => S4313
    );
notg_4772: ENTITY WORK.notg
    PORT MAP (
        in1 => S4313,
        out1 => S4314
    );
nor_n_4773: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4314,
        in1(1) => S5907,
        out1 => S4315
    );
nand_n_4774: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4313,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S4316
    );
nor_n_4775: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4313,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S4317
    );
nor_n_4776: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4313,
        in1(1) => S5907,
        out1 => S4318
    );
nor_n_4777: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4314,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S4319
    );
nor_n_4778: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4317,
        in1(1) => S4315,
        out1 => S4320
    );
notg_4779: ENTITY WORK.notg
    PORT MAP (
        in1 => S4320,
        out1 => S4321
    );
nand_n_4780: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_3,
        in1(1) => S5157,
        out1 => S4323
    );
nand_n_4781: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4288,
        in1(1) => new_controller_fib_3,
        out1 => S4324
    );
nand_n_4782: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4324,
        in1(1) => S4323,
        out1 => S4325
    );
nand_n_4783: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4325,
        in1(1) => S4280,
        out1 => S4326
    );
nand_n_4784: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4294,
        in1(1) => S249,
        out1 => S4327
    );
nand_n_4785: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4327,
        in1(1) => S4326,
        out1 => S4328
    );
notg_4786: ENTITY WORK.notg
    PORT MAP (
        in1 => S4328,
        out1 => S4329
    );
nor_n_4787: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4329,
        in1(1) => S5947,
        out1 => S4330
    );
nand_n_4788: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4328,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S4331
    );
nor_n_4789: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4328,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S4332
    );
notg_4790: ENTITY WORK.notg
    PORT MAP (
        in1 => S4332,
        out1 => S4334
    );
nor_n_4791: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4328,
        in1(1) => S5947,
        out1 => S4335
    );
nor_n_4792: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4329,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S4336
    );
nor_n_4793: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4332,
        in1(1) => S4330,
        out1 => S4337
    );
nand_n_4794: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4334,
        in1(1) => S4331,
        out1 => S4338
    );
nand_n_4795: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_1,
        in1(1) => S5157,
        out1 => S4339
    );
nand_n_4796: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4288,
        in1(1) => new_controller_fib_1,
        out1 => S4340
    );
nand_n_4797: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4340,
        in1(1) => S4339,
        out1 => S4341
    );
nand_n_4798: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4341,
        in1(1) => S4280,
        out1 => S4342
    );
nand_n_4799: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4294,
        in1(1) => S265,
        out1 => S4343
    );
nand_n_4800: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4343,
        in1(1) => S4342,
        out1 => S4345
    );
notg_4801: ENTITY WORK.notg
    PORT MAP (
        in1 => S4345,
        out1 => S4346
    );
nor_n_4802: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4345,
        in1(1) => S5966,
        out1 => S4347
    );
nor_n_4803: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4346,
        in1(1) => S5966,
        out1 => S4348
    );
nand_n_4804: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4345,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S4349
    );
nor_n_4805: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4345,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S4350
    );
notg_4806: ENTITY WORK.notg
    PORT MAP (
        in1 => S4350,
        out1 => S4351
    );
nand_n_4807: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4351,
        in1(1) => S4349,
        out1 => S4352
    );
nor_n_4808: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4350,
        in1(1) => S4348,
        out1 => S4353
    );
nand_n_4809: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_addsubunit_in1_0,
        in1(1) => S5157,
        out1 => S4354
    );
nand_n_4810: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4288,
        in1(1) => new_controller_fib_0,
        out1 => S4356
    );
nand_n_4811: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4356,
        in1(1) => S4354,
        out1 => S4357
    );
nand_n_4812: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4357,
        in1(1) => S4280,
        out1 => S4358
    );
notg_4813: ENTITY WORK.notg
    PORT MAP (
        in1 => S4358,
        out1 => S4359
    );
nor_n_4814: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4293,
        in1(1) => S270,
        out1 => S4360
    );
nand_n_4815: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4294,
        in1(1) => S271,
        out1 => S4361
    );
nor_n_4816: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4360,
        in1(1) => S4359,
        out1 => S4362
    );
nand_n_4817: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4361,
        in1(1) => S4358,
        out1 => S4363
    );
nor_n_4818: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4362,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S4364
    );
nor_n_4819: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4364,
        in1(1) => S4353,
        out1 => S4365
    );
nor_n_4820: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5926,
        in1(1) => S5168,
        out1 => S4367
    );
nand_n_4821: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4286,
        in1(1) => new_controller_234_B_0,
        out1 => S4368
    );
nand_n_4822: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4368,
        in1(1) => S4307,
        out1 => S4369
    );
nor_n_4823: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4369,
        in1(1) => S4367,
        out1 => S4370
    );
nor_n_4824: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4370,
        in1(1) => S4279,
        out1 => S4371
    );
nor_n_4825: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4293,
        in1(1) => S208,
        out1 => S4372
    );
nor_n_4826: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4372,
        in1(1) => S4371,
        out1 => S4373
    );
notg_4827: ENTITY WORK.notg
    PORT MAP (
        in1 => S4373,
        out1 => S4374
    );
nor_n_4828: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4374,
        in1(1) => S5926,
        out1 => S4375
    );
nor_n_4829: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4373,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S4376
    );
nor_n_4830: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4376,
        in1(1) => S4375,
        out1 => S4378
    );
notg_4831: ENTITY WORK.notg
    PORT MAP (
        in1 => S4378,
        out1 => S4379
    );
nor_n_4832: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4363,
        in1(1) => S5975,
        out1 => S4380
    );
nor_n_4833: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4285,
        in1(1) => new_controller_fib_0,
        out1 => S4381
    );
nor_n_4834: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4285,
        in1(1) => S5157,
        out1 => S4382
    );
nor_n_4835: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4382,
        in1(1) => S3062,
        out1 => S4383
    );
nor_n_4836: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4383,
        in1(1) => S5157,
        out1 => S4384
    );
nor_n_4837: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4384,
        in1(1) => S4381,
        out1 => S4385
    );
notg_4838: ENTITY WORK.notg
    PORT MAP (
        in1 => S4385,
        out1 => S4386
    );
nor_n_4839: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4385,
        in1(1) => S4306,
        out1 => S4387
    );
nand_n_4840: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4386,
        in1(1) => S4307,
        out1 => S4389
    );
nor_n_4841: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4387,
        in1(1) => S4279,
        out1 => S4390
    );
nand_n_4842: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4389,
        in1(1) => S4280,
        out1 => S4391
    );
nand_n_4843: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4294,
        in1(1) => new_datapath_multdivunit_1697_B_15,
        out1 => S4392
    );
notg_4844: ENTITY WORK.notg
    PORT MAP (
        in1 => S4392,
        out1 => S4393
    );
nor_n_4845: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4393,
        in1(1) => S4390,
        out1 => S4394
    );
notg_4846: ENTITY WORK.notg
    PORT MAP (
        in1 => S4394,
        out1 => S4395
    );
nand_n_4847: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4394,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S4396
    );
notg_4848: ENTITY WORK.notg
    PORT MAP (
        in1 => S4396,
        out1 => S4397
    );
nor_n_4849: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4394,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S4398
    );
nand_n_4850: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4395,
        in1(1) => S3401,
        out1 => S4400
    );
nor_n_4851: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4398,
        in1(1) => S4397,
        out1 => S4401
    );
nand_n_4852: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4294,
        in1(1) => new_datapath_multdivunit_1697_B_14,
        out1 => S4402
    );
nand_n_4853: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4402,
        in1(1) => S4391,
        out1 => S4403
    );
notg_4854: ENTITY WORK.notg
    PORT MAP (
        in1 => S4403,
        out1 => S4404
    );
nor_n_4855: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4403,
        in1(1) => S3390,
        out1 => S4405
    );
nand_n_4856: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4404,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S4406
    );
nor_n_4857: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4404,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S4407
    );
nor_n_4858: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4404,
        in1(1) => S3390,
        out1 => S4408
    );
nor_n_4859: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4407,
        in1(1) => S4405,
        out1 => S4409
    );
nand_n_4860: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4409,
        in1(1) => S4401,
        out1 => S4411
    );
nand_n_4861: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4294,
        in1(1) => new_datapath_multdivunit_1697_B_13,
        out1 => S4412
    );
nand_n_4862: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4412,
        in1(1) => S4391,
        out1 => S4413
    );
notg_4863: ENTITY WORK.notg
    PORT MAP (
        in1 => S4413,
        out1 => S4414
    );
nor_n_4864: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4413,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S4415
    );
nor_n_4865: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4414,
        in1(1) => S3379,
        out1 => S4416
    );
nor_n_4866: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4416,
        in1(1) => S4415,
        out1 => S4417
    );
notg_4867: ENTITY WORK.notg
    PORT MAP (
        in1 => S4417,
        out1 => S4418
    );
nand_n_4868: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4294,
        in1(1) => new_datapath_multdivunit_1697_B_12,
        out1 => S4419
    );
notg_4869: ENTITY WORK.notg
    PORT MAP (
        in1 => S4419,
        out1 => S4420
    );
nor_n_4870: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4420,
        in1(1) => S4390,
        out1 => S4422
    );
nand_n_4871: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4419,
        in1(1) => S4391,
        out1 => S4423
    );
nor_n_4872: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4422,
        in1(1) => S3368,
        out1 => S4424
    );
nor_n_4873: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4423,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S4425
    );
nand_n_4874: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4422,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S4426
    );
nor_n_4875: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4425,
        in1(1) => S4424,
        out1 => S4427
    );
nor_n_4876: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4427,
        in1(1) => S4417,
        out1 => S4428
    );
notg_4877: ENTITY WORK.notg
    PORT MAP (
        in1 => S4428,
        out1 => S4429
    );
nor_n_4878: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4429,
        in1(1) => S4411,
        out1 => S4430
    );
nand_n_4879: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4294,
        in1(1) => new_datapath_multdivunit_1697_B_10,
        out1 => S4431
    );
nand_n_4880: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4431,
        in1(1) => S4391,
        out1 => S4433
    );
nor_n_4881: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4433,
        in1(1) => S3346,
        out1 => S4434
    );
nand_n_4882: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4433,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S4435
    );
notg_4883: ENTITY WORK.notg
    PORT MAP (
        in1 => S4435,
        out1 => S4436
    );
nor_n_4884: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4433,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S4437
    );
nor_n_4885: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4437,
        in1(1) => S4436,
        out1 => S4438
    );
nand_n_4886: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4294,
        in1(1) => new_datapath_multdivunit_1697_B_8,
        out1 => S4439
    );
nand_n_4887: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4439,
        in1(1) => S4391,
        out1 => S4440
    );
notg_4888: ENTITY WORK.notg
    PORT MAP (
        in1 => S4440,
        out1 => S4441
    );
nand_n_4889: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4440,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S4442
    );
notg_4890: ENTITY WORK.notg
    PORT MAP (
        in1 => S4442,
        out1 => S4444
    );
nor_n_4891: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4440,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S4445
    );
nand_n_4892: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4441,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S4446
    );
nor_n_4893: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4445,
        in1(1) => S4444,
        out1 => S4447
    );
notg_4894: ENTITY WORK.notg
    PORT MAP (
        in1 => S4447,
        out1 => S4448
    );
nand_n_4895: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4294,
        in1(1) => new_datapath_multdivunit_1697_B_9,
        out1 => S4449
    );
nand_n_4896: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4449,
        in1(1) => S4391,
        out1 => S4450
    );
notg_4897: ENTITY WORK.notg
    PORT MAP (
        in1 => S4450,
        out1 => S4451
    );
nor_n_4898: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4450,
        in1(1) => S3336,
        out1 => S4452
    );
nor_n_4899: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4451,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S4453
    );
nor_n_4900: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4453,
        in1(1) => S4452,
        out1 => S4455
    );
notg_4901: ENTITY WORK.notg
    PORT MAP (
        in1 => S4455,
        out1 => S4456
    );
nand_n_4902: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4455,
        in1(1) => S4448,
        out1 => S4457
    );
nand_n_4903: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4294,
        in1(1) => new_datapath_multdivunit_1697_B_11,
        out1 => S4458
    );
notg_4904: ENTITY WORK.notg
    PORT MAP (
        in1 => S4458,
        out1 => S4459
    );
nor_n_4905: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4459,
        in1(1) => S4390,
        out1 => S4460
    );
nand_n_4906: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4458,
        in1(1) => S4391,
        out1 => S4461
    );
nor_n_4907: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4460,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S4462
    );
nor_n_4908: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4461,
        in1(1) => S3357,
        out1 => S4463
    );
nor_n_4909: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4460,
        in1(1) => S3357,
        out1 => S4464
    );
nor_n_4910: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4461,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S4466
    );
nor_n_4911: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4466,
        in1(1) => S4464,
        out1 => S4467
    );
nor_n_4912: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5916,
        in1(1) => S5168,
        out1 => S4468
    );
nand_n_4913: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4286,
        in1(1) => new_controller_opcode_2,
        out1 => S4469
    );
nand_n_4914: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4469,
        in1(1) => S4307,
        out1 => S4470
    );
nor_n_4915: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4470,
        in1(1) => S4468,
        out1 => S4471
    );
notg_4916: ENTITY WORK.notg
    PORT MAP (
        in1 => S4471,
        out1 => S4472
    );
nand_n_4917: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4472,
        in1(1) => S4280,
        out1 => S4473
    );
nand_n_4918: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4294,
        in1(1) => S203,
        out1 => S4474
    );
nand_n_4919: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4474,
        in1(1) => S4473,
        out1 => S4475
    );
notg_4920: ENTITY WORK.notg
    PORT MAP (
        in1 => S4475,
        out1 => S4477
    );
nor_n_4921: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4475,
        in1(1) => S5916,
        out1 => S4478
    );
nor_n_4922: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4477,
        in1(1) => S5916,
        out1 => S4479
    );
nand_n_4923: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4475,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S4480
    );
nor_n_4924: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4475,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S4481
    );
nor_n_4925: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4481,
        in1(1) => S4479,
        out1 => S4482
    );
notg_4926: ENTITY WORK.notg
    PORT MAP (
        in1 => S4482,
        out1 => S4483
    );
nor_n_4927: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5936,
        in1(1) => S5168,
        out1 => S4484
    );
nand_n_4928: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4288,
        in1(1) => new_controller_fib_4,
        out1 => S4485
    );
notg_4929: ENTITY WORK.notg
    PORT MAP (
        in1 => S4485,
        out1 => S4486
    );
nor_n_4930: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4486,
        in1(1) => S4484,
        out1 => S4488
    );
notg_4931: ENTITY WORK.notg
    PORT MAP (
        in1 => S4488,
        out1 => S4489
    );
nor_n_4932: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4488,
        in1(1) => S4279,
        out1 => S4490
    );
nand_n_4933: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4489,
        in1(1) => S4280,
        out1 => S4491
    );
nor_n_4934: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4293,
        in1(1) => S240,
        out1 => S4492
    );
nand_n_4935: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4294,
        in1(1) => S241,
        out1 => S4493
    );
nor_n_4936: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4492,
        in1(1) => S4490,
        out1 => S4494
    );
nand_n_4937: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4493,
        in1(1) => S4491,
        out1 => S4495
    );
nor_n_4938: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4494,
        in1(1) => S5936,
        out1 => S4496
    );
notg_4939: ENTITY WORK.notg
    PORT MAP (
        in1 => S4496,
        out1 => S4497
    );
nor_n_4940: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4495,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S4499
    );
nand_n_4941: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4494,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S4500
    );
nor_n_4942: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4499,
        in1(1) => S4496,
        out1 => S4501
    );
notg_4943: ENTITY WORK.notg
    PORT MAP (
        in1 => S4501,
        out1 => S4502
    );
nand_n_4944: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4363,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S4503
    );
nor_n_4945: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4380,
        in1(1) => S4364,
        out1 => S4504
    );
notg_4946: ENTITY WORK.notg
    PORT MAP (
        in1 => S4504,
        out1 => S4505
    );
nor_n_4947: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4501,
        in1(1) => S4302,
        out1 => S4506
    );
nor_n_4948: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4482,
        in1(1) => S4320,
        out1 => S4507
    );
nand_n_4949: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4506,
        in1(1) => S4378,
        out1 => S4508
    );
nor_n_4950: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4337,
        in1(1) => S4274,
        out1 => S4510
    );
nor_n_4951: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4467,
        in1(1) => S4438,
        out1 => S4511
    );
nand_n_4952: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4511,
        in1(1) => S4430,
        out1 => S4512
    );
nor_n_4953: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4512,
        in1(1) => S4457,
        out1 => S4513
    );
nand_n_4954: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4513,
        in1(1) => S4504,
        out1 => S4514
    );
nor_n_4955: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4514,
        in1(1) => S4353,
        out1 => S4515
    );
nand_n_4956: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4515,
        in1(1) => S4510,
        out1 => S4516
    );
nor_n_4957: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4516,
        in1(1) => S4508,
        out1 => S4517
    );
nand_n_4958: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4517,
        in1(1) => S4507,
        out1 => S4518
    );
nand_n_4959: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4518,
        in1(1) => S4275,
        out1 => S70
    );
nand_n_4960: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4274,
        in1(1) => new_controller_407_B_2,
        out1 => S4520
    );
nor_n_4961: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4365,
        in1(1) => S4347,
        out1 => S4521
    );
nor_n_4962: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4521,
        in1(1) => S4302,
        out1 => S4522
    );
nor_n_4963: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4522,
        in1(1) => S4297,
        out1 => S4523
    );
notg_4964: ENTITY WORK.notg
    PORT MAP (
        in1 => S4523,
        out1 => S4524
    );
nor_n_4965: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4523,
        in1(1) => S4336,
        out1 => S4525
    );
nor_n_4966: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4525,
        in1(1) => S4335,
        out1 => S4526
    );
notg_4967: ENTITY WORK.notg
    PORT MAP (
        in1 => S4526,
        out1 => S4527
    );
nand_n_4968: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4527,
        in1(1) => S4502,
        out1 => S4528
    );
nand_n_4969: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4528,
        in1(1) => S4500,
        out1 => S4529
    );
notg_4970: ENTITY WORK.notg
    PORT MAP (
        in1 => S4529,
        out1 => S4531
    );
nor_n_4971: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4531,
        in1(1) => S4376,
        out1 => S4532
    );
nor_n_4972: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4532,
        in1(1) => S4375,
        out1 => S4533
    );
nor_n_4973: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4533,
        in1(1) => S4482,
        out1 => S4534
    );
nor_n_4974: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4534,
        in1(1) => S4478,
        out1 => S4535
    );
notg_4975: ENTITY WORK.notg
    PORT MAP (
        in1 => S4535,
        out1 => S4536
    );
nor_n_4976: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4535,
        in1(1) => S4319,
        out1 => S4537
    );
nor_n_4977: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4537,
        in1(1) => S4318,
        out1 => S4538
    );
nor_n_4978: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4538,
        in1(1) => S4447,
        out1 => S4539
    );
notg_4979: ENTITY WORK.notg
    PORT MAP (
        in1 => S4539,
        out1 => S4540
    );
nand_n_4980: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4540,
        in1(1) => S4446,
        out1 => S4542
    );
notg_4981: ENTITY WORK.notg
    PORT MAP (
        in1 => S4542,
        out1 => S4543
    );
nor_n_4982: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4543,
        in1(1) => S4453,
        out1 => S4544
    );
nor_n_4983: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4544,
        in1(1) => S4452,
        out1 => S4545
    );
nor_n_4984: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4545,
        in1(1) => S4438,
        out1 => S4546
    );
nor_n_4985: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4546,
        in1(1) => S4434,
        out1 => S4547
    );
nor_n_4986: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4547,
        in1(1) => S4462,
        out1 => S4548
    );
nor_n_4987: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4548,
        in1(1) => S4463,
        out1 => S4549
    );
notg_4988: ENTITY WORK.notg
    PORT MAP (
        in1 => S4549,
        out1 => S4550
    );
nand_n_4989: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4550,
        in1(1) => S4430,
        out1 => S4551
    );
nor_n_4990: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4413,
        in1(1) => S3379,
        out1 => S4553
    );
nand_n_4991: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4414,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S4554
    );
nor_n_4992: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4426,
        in1(1) => S4417,
        out1 => S4555
    );
nor_n_4993: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4555,
        in1(1) => S4553,
        out1 => S4556
    );
nor_n_4994: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4556,
        in1(1) => S4411,
        out1 => S4557
    );
nand_n_4995: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4406,
        in1(1) => S4396,
        out1 => S4558
    );
nand_n_4996: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4558,
        in1(1) => S4400,
        out1 => S4559
    );
nand_n_4997: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4559,
        in1(1) => S4273,
        out1 => S4560
    );
nor_n_4998: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4560,
        in1(1) => S4557,
        out1 => S4561
    );
nand_n_4999: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4561,
        in1(1) => S4551,
        out1 => S4562
    );
nand_n_5000: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4562,
        in1(1) => S4520,
        out1 => S71
    );
nand_n_5001: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6091,
        in1(1) => new_datapath_adr_outreg_0,
        out1 => S4564
    );
nand_n_5002: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6090,
        in1(1) => S5977,
        out1 => S4565
    );
nand_n_5003: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4565,
        in1(1) => S4564,
        out1 => S73
    );
nand_n_5004: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6091,
        in1(1) => new_datapath_adr_outreg_1,
        out1 => S4566
    );
nand_n_5005: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6090,
        in1(1) => S5968,
        out1 => S4567
    );
nand_n_5006: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4567,
        in1(1) => S4566,
        out1 => S74
    );
nand_n_5007: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6091,
        in1(1) => new_datapath_adr_outreg_2,
        out1 => S4568
    );
nand_n_5008: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6090,
        in1(1) => S5959,
        out1 => S4569
    );
nand_n_5009: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4569,
        in1(1) => S4568,
        out1 => S75
    );
nand_n_5010: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6091,
        in1(1) => new_datapath_adr_outreg_3,
        out1 => S4571
    );
nand_n_5011: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6090,
        in1(1) => S5949,
        out1 => S4572
    );
nand_n_5012: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4572,
        in1(1) => S4571,
        out1 => S76
    );
nand_n_5013: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6091,
        in1(1) => new_datapath_adr_outreg_4,
        out1 => S4573
    );
nand_n_5014: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6090,
        in1(1) => S5938,
        out1 => S4574
    );
nand_n_5015: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4574,
        in1(1) => S4573,
        out1 => S77
    );
nand_n_5016: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6091,
        in1(1) => new_datapath_adr_outreg_5,
        out1 => S4575
    );
nand_n_5017: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6090,
        in1(1) => S5928,
        out1 => S4576
    );
nand_n_5018: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4576,
        in1(1) => S4575,
        out1 => S78
    );
nand_n_5019: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6091,
        in1(1) => new_datapath_adr_outreg_6,
        out1 => S4577
    );
nand_n_5020: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6090,
        in1(1) => S5918,
        out1 => S4579
    );
nand_n_5021: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4579,
        in1(1) => S4577,
        out1 => S79
    );
nand_n_5022: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6091,
        in1(1) => new_datapath_adr_outreg_7,
        out1 => S4580
    );
nand_n_5023: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6090,
        in1(1) => S5909,
        out1 => S4581
    );
nand_n_5024: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4581,
        in1(1) => S4580,
        out1 => S80
    );
nand_n_5025: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6091,
        in1(1) => new_datapath_adr_outreg_8,
        out1 => S4582
    );
nand_n_5026: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6090,
        in1(1) => S4975,
        out1 => S4583
    );
nand_n_5027: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4583,
        in1(1) => S4582,
        out1 => S81
    );
nand_n_5028: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6091,
        in1(1) => new_datapath_adr_outreg_9,
        out1 => S4584
    );
nand_n_5029: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6090,
        in1(1) => S4922,
        out1 => S4585
    );
nand_n_5030: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4585,
        in1(1) => S4584,
        out1 => S82
    );
nand_n_5031: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6091,
        in1(1) => new_datapath_adr_outreg_10,
        out1 => S4587
    );
nand_n_5032: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6090,
        in1(1) => S4857,
        out1 => S4588
    );
nand_n_5033: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4588,
        in1(1) => S4587,
        out1 => S83
    );
nand_n_5034: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6091,
        in1(1) => new_datapath_adr_outreg_11,
        out1 => S4589
    );
nand_n_5035: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6090,
        in1(1) => S4804,
        out1 => S4590
    );
nand_n_5036: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4590,
        in1(1) => S4589,
        out1 => S84
    );
nand_n_5037: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6091,
        in1(1) => new_datapath_adr_outreg_12,
        out1 => S4591
    );
nand_n_5038: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6090,
        in1(1) => S4740,
        out1 => S4592
    );
nand_n_5039: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4592,
        in1(1) => S4591,
        out1 => S85
    );
nand_n_5040: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6091,
        in1(1) => new_datapath_adr_outreg_13,
        out1 => S4594
    );
nand_n_5041: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6090,
        in1(1) => S4686,
        out1 => S4595
    );
nand_n_5042: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4595,
        in1(1) => S4594,
        out1 => S86
    );
nand_n_5043: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6091,
        in1(1) => new_datapath_adr_outreg_14,
        out1 => S4596
    );
nand_n_5044: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6090,
        in1(1) => S4621,
        out1 => S4597
    );
nand_n_5045: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4597,
        in1(1) => S4596,
        out1 => S87
    );
nand_n_5046: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5136,
        in1(1) => S4089,
        out1 => S4598
    );
notg_5047: ENTITY WORK.notg
    PORT MAP (
        in1 => S4598,
        out1 => S4599
    );
nor_n_5048: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5451,
        in1(1) => S5239,
        out1 => S4600
    );
notg_5049: ENTITY WORK.notg
    PORT MAP (
        in1 => S4600,
        out1 => S4601
    );
nand_n_5050: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4598,
        in1(1) => S3870,
        out1 => S4603
    );
nand_n_5051: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4600,
        in1(1) => S5663,
        out1 => S4604
    );
nor_n_5052: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4604,
        in1(1) => S4603,
        out1 => S4605
    );
nand_n_5053: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5483,
        in1(1) => S5311,
        out1 => S4606
    );
nor_n_5054: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S170,
        in1(1) => S3947,
        out1 => S4607
    );
nor_n_5055: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4607,
        in1(1) => S4606,
        out1 => S4608
    );
nand_n_5056: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4608,
        in1(1) => S4605,
        out1 => S4609
    );
nand_n_5057: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4609,
        in1(1) => S3761,
        out1 => S4610
    );
nor_n_5058: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4166,
        in1(1) => S3740,
        out1 => S4611
    );
nor_n_5059: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4611,
        in1(1) => S4122,
        out1 => S4612
    );
nand_n_5060: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4612,
        in1(1) => S4610,
        out1 => new_controller_1133_Y
    );
nor_n_5061: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => S6086,
        out1 => S4614
    );
notg_5062: ENTITY WORK.notg
    PORT MAP (
        in1 => S4614,
        out1 => new_controller_1423_Y_0
    );
nand_n_5063: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4166,
        in1(1) => S3708,
        out1 => S4615
    );
nand_n_5064: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6091,
        in1(1) => S5611,
        out1 => S4616
    );
nor_n_5065: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4616,
        in1(1) => S6086,
        out1 => S4617
    );
nand_n_5066: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4617,
        in1(1) => S4615,
        out1 => new_controller_1423_Y_1
    );
nor_n_5067: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5280,
        in1(1) => S3620,
        out1 => S4618
    );
nand_n_5068: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5271,
        in1(1) => S3609,
        out1 => S4619
    );
nor_n_5069: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4618,
        in1(1) => S5255,
        out1 => S4620
    );
nand_n_5070: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4619,
        in1(1) => S5262,
        out1 => S4622
    );
nor_n_5071: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4620,
        in1(1) => S3771,
        out1 => S4623
    );
nand_n_5072: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4622,
        in1(1) => S3761,
        out1 => S4624
    );
nor_n_5073: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5558,
        in1(1) => S5280,
        out1 => S4625
    );
nand_n_5074: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5568,
        in1(1) => S5271,
        out1 => S4626
    );
nand_n_5075: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4626,
        in1(1) => S4624,
        out1 => S4627
    );
nand_n_5076: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4627,
        in1(1) => S4505,
        out1 => S4628
    );
nor_n_5077: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4600,
        in1(1) => S3771,
        out1 => S4629
    );
nand_n_5078: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4601,
        in1(1) => S3761,
        out1 => S4630
    );
nor_n_5079: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4630,
        in1(1) => S4503,
        out1 => S4631
    );
nor_n_5080: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4598,
        in1(1) => S3771,
        out1 => S4633
    );
nand_n_5081: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4599,
        in1(1) => S3761,
        out1 => S4634
    );
nand_n_5082: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4633,
        in1(1) => S4357,
        out1 => S4635
    );
nor_n_5083: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5975,
        in1(1) => new_controller_fib_4,
        out1 => S4636
    );
nor_n_5084: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4578,
        in1(1) => S4269,
        out1 => S4637
    );
nand_n_5085: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4570,
        in1(1) => S4278,
        out1 => S4638
    );
nand_n_5086: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4637,
        in1(1) => new_controller_fib_4,
        out1 => S4639
    );
notg_5087: ENTITY WORK.notg
    PORT MAP (
        in1 => S4639,
        out1 => S4640
    );
nand_n_5088: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4640,
        in1(1) => S5975,
        out1 => S4641
    );
notg_5089: ENTITY WORK.notg
    PORT MAP (
        in1 => S4641,
        out1 => S4642
    );
nand_n_5090: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4641,
        in1(1) => S4637,
        out1 => S4644
    );
nor_n_5091: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4644,
        in1(1) => S4636,
        out1 => S4645
    );
nand_n_5092: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S241,
        in1(1) => S5683,
        out1 => S4646
    );
nand_n_5093: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5115,
        in1(1) => new_controller_fib_4,
        out1 => S4647
    );
nand_n_5094: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4647,
        in1(1) => S4646,
        out1 => S4648
    );
notg_5095: ENTITY WORK.notg
    PORT MAP (
        in1 => S4648,
        out1 => S4649
    );
nor_n_5096: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5632,
        in1(1) => S3771,
        out1 => S4650
    );
nor_n_5097: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5125,
        in1(1) => S3040,
        out1 => S4651
    );
nor_n_5098: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4651,
        in1(1) => S4650,
        out1 => S4652
    );
notg_5099: ENTITY WORK.notg
    PORT MAP (
        in1 => S4652,
        out1 => S4653
    );
nor_n_5100: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5653,
        in1(1) => S3771,
        out1 => S4655
    );
nor_n_5101: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5125,
        in1(1) => new_controller_234_B_0,
        out1 => S4656
    );
nor_n_5102: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4656,
        in1(1) => S4655,
        out1 => S4657
    );
nand_n_5103: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4657,
        in1(1) => S4652,
        out1 => S4658
    );
notg_5104: ENTITY WORK.notg
    PORT MAP (
        in1 => S4658,
        out1 => S4659
    );
nor_n_5105: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4659,
        in1(1) => S4648,
        out1 => S4660
    );
nand_n_5106: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4658,
        in1(1) => S4649,
        out1 => S4661
    );
nand_n_5107: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4660,
        in1(1) => new_datapath_shiftunit_1961_A,
        out1 => S4662
    );
nand_n_5108: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4648,
        in1(1) => new_datapath_shiftunit_2265_A,
        out1 => S4663
    );
notg_5109: ENTITY WORK.notg
    PORT MAP (
        in1 => S4663,
        out1 => S4664
    );
nand_n_5110: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6215,
        in1(1) => new_datapath_databusin_0,
        out1 => S4666
    );
nand_n_5111: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => new_datapath_multdivunit_outmdu1_0,
        out1 => S4667
    );
nand_n_5112: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4144,
        in1(1) => new_datapath_multdivunit_outmdu2_0,
        out1 => S4668
    );
nor_n_5113: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S170,
        in1(1) => S4261,
        out1 => S4669
    );
nand_n_5114: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4607,
        in1(1) => S3761,
        out1 => S4670
    );
nor_n_5115: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4670,
        in1(1) => new_datapath_muxmem_in2_0,
        out1 => S4671
    );
nand_n_5116: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4668,
        in1(1) => S4667,
        out1 => S4672
    );
nor_n_5117: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4672,
        in1(1) => S4671,
        out1 => S4673
    );
nand_n_5118: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4673,
        in1(1) => S4666,
        out1 => S4674
    );
nor_n_5119: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4674,
        in1(1) => S4664,
        out1 => S4675
    );
nand_n_5120: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4675,
        in1(1) => S4662,
        out1 => S4677
    );
nor_n_5121: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4677,
        in1(1) => S4645,
        out1 => S4678
    );
nand_n_5122: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4678,
        in1(1) => S4635,
        out1 => S4679
    );
nor_n_5123: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4679,
        in1(1) => S4631,
        out1 => S4680
    );
nand_n_5124: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4680,
        in1(1) => S4628,
        out1 => new_datapath_indatatrf_0
    );
nand_n_5125: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4364,
        in1(1) => S4353,
        out1 => S4681
    );
nor_n_5126: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4624,
        in1(1) => S4365,
        out1 => S4682
    );
nand_n_5127: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4682,
        in1(1) => S4681,
        out1 => S4683
    );
nor_n_5128: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4503,
        in1(1) => S4352,
        out1 => S4684
    );
notg_5129: ENTITY WORK.notg
    PORT MAP (
        in1 => S4684,
        out1 => S4685
    );
nand_n_5130: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4503,
        in1(1) => S4352,
        out1 => S4687
    );
nand_n_5131: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4687,
        in1(1) => S4625,
        out1 => S4688
    );
nor_n_5132: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4688,
        in1(1) => S4684,
        out1 => S4689
    );
nand_n_5133: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4629,
        in1(1) => S4348,
        out1 => S4690
    );
nor_n_5134: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4644,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S4691
    );
nand_n_5135: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4633,
        in1(1) => S4341,
        out1 => S4692
    );
nor_n_5136: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4641,
        in1(1) => S5966,
        out1 => S4693
    );
nand_n_5137: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4660,
        in1(1) => new_datapath_shiftunit_1979_A,
        out1 => S4694
    );
nand_n_5138: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4648,
        in1(1) => new_datapath_shiftunit_2283_A,
        out1 => S4695
    );
nand_n_5139: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4144,
        in1(1) => new_datapath_multdivunit_outmdu2_1,
        out1 => S4696
    );
nand_n_5140: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => new_datapath_multdivunit_outmdu1_1,
        out1 => S4698
    );
nand_n_5141: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4698,
        in1(1) => S4696,
        out1 => S4699
    );
nand_n_5142: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6215,
        in1(1) => new_datapath_databusin_1,
        out1 => S4700
    );
nand_n_5143: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4669,
        in1(1) => S6110,
        out1 => S4701
    );
nand_n_5144: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4701,
        in1(1) => S4700,
        out1 => S4702
    );
nor_n_5145: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4702,
        in1(1) => S4699,
        out1 => S4703
    );
nand_n_5146: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4703,
        in1(1) => S4695,
        out1 => S4704
    );
notg_5147: ENTITY WORK.notg
    PORT MAP (
        in1 => S4704,
        out1 => S4705
    );
nand_n_5148: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4705,
        in1(1) => S4694,
        out1 => S4706
    );
nor_n_5149: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4706,
        in1(1) => S4693,
        out1 => S4707
    );
nand_n_5150: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4707,
        in1(1) => S4692,
        out1 => S4709
    );
nor_n_5151: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4641,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S4710
    );
nand_n_5152: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4642,
        in1(1) => S5966,
        out1 => S4711
    );
nor_n_5153: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4709,
        in1(1) => S4691,
        out1 => S4712
    );
nand_n_5154: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4712,
        in1(1) => S4690,
        out1 => S4713
    );
nor_n_5155: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4713,
        in1(1) => S4689,
        out1 => S4714
    );
nand_n_5156: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4714,
        in1(1) => S4683,
        out1 => new_datapath_indatatrf_1
    );
nand_n_5157: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4685,
        in1(1) => S4349,
        out1 => S4715
    );
nand_n_5158: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4715,
        in1(1) => S4302,
        out1 => S4716
    );
nor_n_5159: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4715,
        in1(1) => S4302,
        out1 => S4717
    );
nand_n_5160: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4716,
        in1(1) => S4625,
        out1 => S4719
    );
nor_n_5161: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4719,
        in1(1) => S4717,
        out1 => S4720
    );
nand_n_5162: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4521,
        in1(1) => S4302,
        out1 => S4721
    );
nor_n_5163: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4624,
        in1(1) => S4522,
        out1 => S4722
    );
nand_n_5164: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4722,
        in1(1) => S4721,
        out1 => S4723
    );
nand_n_5165: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4629,
        in1(1) => S4299,
        out1 => S4724
    );
nand_n_5166: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4633,
        in1(1) => S4291,
        out1 => S4725
    );
nor_n_5167: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4661,
        in1(1) => S3489,
        out1 => S4726
    );
nand_n_5168: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4648,
        in1(1) => new_datapath_shiftunit_2301_A,
        out1 => S4727
    );
nand_n_5169: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4669,
        in1(1) => S6124,
        out1 => S4728
    );
nand_n_5170: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => new_datapath_multdivunit_outmdu1_2,
        out1 => S4730
    );
nand_n_5171: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4730,
        in1(1) => S4728,
        out1 => S4731
    );
nand_n_5172: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4144,
        in1(1) => new_datapath_multdivunit_outmdu2_2,
        out1 => S4732
    );
nand_n_5173: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6215,
        in1(1) => new_datapath_databusin_2,
        out1 => S4733
    );
nand_n_5174: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4733,
        in1(1) => S4732,
        out1 => S4734
    );
nor_n_5175: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4734,
        in1(1) => S4731,
        out1 => S4735
    );
nand_n_5176: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4735,
        in1(1) => S4727,
        out1 => S4736
    );
nor_n_5177: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4736,
        in1(1) => S4726,
        out1 => S4737
    );
nand_n_5178: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4737,
        in1(1) => S4725,
        out1 => S4738
    );
nor_n_5179: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4710,
        in1(1) => S5957,
        out1 => S4739
    );
nor_n_5180: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4711,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S4741
    );
nand_n_5181: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4710,
        in1(1) => S5957,
        out1 => S4742
    );
nand_n_5182: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4742,
        in1(1) => S4637,
        out1 => S4743
    );
nor_n_5183: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4743,
        in1(1) => S4739,
        out1 => S4744
    );
nor_n_5184: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4744,
        in1(1) => S4738,
        out1 => S4745
    );
nand_n_5185: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4745,
        in1(1) => S4724,
        out1 => S4746
    );
nor_n_5186: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4746,
        in1(1) => S4720,
        out1 => S4747
    );
nand_n_5187: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4747,
        in1(1) => S4723,
        out1 => new_datapath_indatatrf_2
    );
nor_n_5188: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4523,
        in1(1) => S4338,
        out1 => S4748
    );
nor_n_5189: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4524,
        in1(1) => S4337,
        out1 => S4749
    );
nor_n_5190: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4749,
        in1(1) => S4748,
        out1 => S4751
    );
nor_n_5191: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4751,
        in1(1) => S4624,
        out1 => S4752
    );
nand_n_5192: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4716,
        in1(1) => S4298,
        out1 => S4753
    );
notg_5193: ENTITY WORK.notg
    PORT MAP (
        in1 => S4753,
        out1 => S4754
    );
nand_n_5194: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4753,
        in1(1) => S4338,
        out1 => S4755
    );
nand_n_5195: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4754,
        in1(1) => S4337,
        out1 => S4756
    );
nand_n_5196: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4756,
        in1(1) => S4755,
        out1 => S4757
    );
nand_n_5197: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4757,
        in1(1) => S4625,
        out1 => S4758
    );
nand_n_5198: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4742,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S4759
    );
nor_n_5199: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4742,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S4760
    );
nand_n_5200: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4741,
        in1(1) => S5947,
        out1 => S4762
    );
nor_n_5201: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4760,
        in1(1) => S4638,
        out1 => S4763
    );
nand_n_5202: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4763,
        in1(1) => S4759,
        out1 => S4764
    );
nor_n_5203: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4630,
        in1(1) => S4331,
        out1 => S4765
    );
nand_n_5204: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4633,
        in1(1) => S4325,
        out1 => S4766
    );
nor_n_5205: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4661,
        in1(1) => S3500,
        out1 => S4767
    );
nand_n_5206: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4648,
        in1(1) => new_datapath_shiftunit_2319_A,
        out1 => S4768
    );
nand_n_5207: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4669,
        in1(1) => S6140,
        out1 => S4769
    );
nand_n_5208: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6215,
        in1(1) => new_datapath_databusin_3,
        out1 => S4770
    );
nand_n_5209: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4770,
        in1(1) => S4769,
        out1 => S4771
    );
nand_n_5210: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => new_datapath_multdivunit_outmdu1_3,
        out1 => S4773
    );
nand_n_5211: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4144,
        in1(1) => new_datapath_multdivunit_outmdu2_3,
        out1 => S4774
    );
nand_n_5212: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4774,
        in1(1) => S4773,
        out1 => S4775
    );
nor_n_5213: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4775,
        in1(1) => S4771,
        out1 => S4776
    );
nand_n_5214: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4776,
        in1(1) => S4768,
        out1 => S4777
    );
nor_n_5215: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4777,
        in1(1) => S4767,
        out1 => S4778
    );
nand_n_5216: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4778,
        in1(1) => S4766,
        out1 => S4779
    );
nor_n_5217: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4779,
        in1(1) => S4765,
        out1 => S4780
    );
nand_n_5218: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4780,
        in1(1) => S4764,
        out1 => S4781
    );
nor_n_5219: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4781,
        in1(1) => S4752,
        out1 => S4782
    );
nand_n_5220: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4782,
        in1(1) => S4758,
        out1 => new_datapath_indatatrf_3
    );
nand_n_5221: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4526,
        in1(1) => S4501,
        out1 => S4784
    );
nand_n_5222: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4784,
        in1(1) => S4528,
        out1 => S4785
    );
nor_n_5223: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4785,
        in1(1) => S4624,
        out1 => S4786
    );
nand_n_5224: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4753,
        in1(1) => S4334,
        out1 => S4787
    );
nand_n_5225: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4787,
        in1(1) => S4331,
        out1 => S4788
    );
nor_n_5226: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4788,
        in1(1) => S4501,
        out1 => S4789
    );
nand_n_5227: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4788,
        in1(1) => S4501,
        out1 => S4790
    );
nor_n_5228: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4789,
        in1(1) => S4626,
        out1 => S4791
    );
nand_n_5229: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4791,
        in1(1) => S4790,
        out1 => S4792
    );
nor_n_5230: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4760,
        in1(1) => S5936,
        out1 => S4794
    );
nor_n_5231: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4762,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S4795
    );
nand_n_5232: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4760,
        in1(1) => S5936,
        out1 => S4796
    );
nand_n_5233: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4796,
        in1(1) => S4637,
        out1 => S4797
    );
nor_n_5234: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4797,
        in1(1) => S4794,
        out1 => S4798
    );
nand_n_5235: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4629,
        in1(1) => S4496,
        out1 => S4799
    );
nor_n_5236: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4634,
        in1(1) => S4488,
        out1 => S4800
    );
nand_n_5237: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4660,
        in1(1) => new_datapath_shiftunit_2033_A,
        out1 => S4801
    );
nand_n_5238: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4648,
        in1(1) => new_datapath_shiftunit_2337_A,
        out1 => S4802
    );
nand_n_5239: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6215,
        in1(1) => new_datapath_databusin_4,
        out1 => S4803
    );
nand_n_5240: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => new_datapath_multdivunit_outmdu1_4,
        out1 => S4805
    );
nand_n_5241: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4144,
        in1(1) => new_datapath_multdivunit_outmdu2_4,
        out1 => S4806
    );
nor_n_5242: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4670,
        in1(1) => S6153,
        out1 => S4807
    );
nand_n_5243: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4806,
        in1(1) => S4805,
        out1 => S4808
    );
nor_n_5244: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4808,
        in1(1) => S4807,
        out1 => S4809
    );
nand_n_5245: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4809,
        in1(1) => S4802,
        out1 => S4810
    );
notg_5246: ENTITY WORK.notg
    PORT MAP (
        in1 => S4810,
        out1 => S4811
    );
nand_n_5247: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4811,
        in1(1) => S4801,
        out1 => S4812
    );
nor_n_5248: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4812,
        in1(1) => S4800,
        out1 => S4813
    );
nand_n_5249: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4813,
        in1(1) => S4799,
        out1 => S4814
    );
nor_n_5250: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4814,
        in1(1) => S4798,
        out1 => S4816
    );
nand_n_5251: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4816,
        in1(1) => S4803,
        out1 => S4817
    );
nor_n_5252: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4817,
        in1(1) => S4786,
        out1 => S4818
    );
nand_n_5253: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4818,
        in1(1) => S4792,
        out1 => new_datapath_indatatrf_4
    );
nor_n_5254: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4529,
        in1(1) => S4378,
        out1 => S4819
    );
nand_n_5255: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4529,
        in1(1) => S4378,
        out1 => S4820
    );
nand_n_5256: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4820,
        in1(1) => S4623,
        out1 => S4821
    );
nor_n_5257: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4821,
        in1(1) => S4819,
        out1 => S4822
    );
nand_n_5258: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4790,
        in1(1) => S4497,
        out1 => S4823
    );
nand_n_5259: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4823,
        in1(1) => S4379,
        out1 => S4824
    );
notg_5260: ENTITY WORK.notg
    PORT MAP (
        in1 => S4824,
        out1 => S4826
    );
nor_n_5261: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4823,
        in1(1) => S4379,
        out1 => S4827
    );
nand_n_5262: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4824,
        in1(1) => S4625,
        out1 => S4828
    );
nor_n_5263: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4828,
        in1(1) => S4827,
        out1 => S4829
    );
nor_n_5264: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4373,
        in1(1) => S5926,
        out1 => S4830
    );
nand_n_5265: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4830,
        in1(1) => S4629,
        out1 => S4831
    );
nor_n_5266: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4634,
        in1(1) => S4370,
        out1 => S4832
    );
nand_n_5267: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4660,
        in1(1) => new_datapath_shiftunit_2051_A,
        out1 => S4833
    );
nand_n_5268: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4648,
        in1(1) => new_datapath_shiftunit_2355_A,
        out1 => S4834
    );
notg_5269: ENTITY WORK.notg
    PORT MAP (
        in1 => S4834,
        out1 => S4835
    );
nor_n_5270: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4670,
        in1(1) => S6167,
        out1 => S4837
    );
nand_n_5271: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4144,
        in1(1) => new_datapath_multdivunit_outmdu2_5,
        out1 => S4838
    );
nand_n_5272: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6215,
        in1(1) => new_datapath_databusin_5,
        out1 => S4839
    );
nand_n_5273: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => new_datapath_multdivunit_outmdu1_5,
        out1 => S4840
    );
nand_n_5274: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4840,
        in1(1) => S4838,
        out1 => S4841
    );
nor_n_5275: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4841,
        in1(1) => S4837,
        out1 => S4842
    );
nand_n_5276: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4842,
        in1(1) => S4839,
        out1 => S4843
    );
nor_n_5277: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4843,
        in1(1) => S4835,
        out1 => S4844
    );
nand_n_5278: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4844,
        in1(1) => S4833,
        out1 => S4845
    );
nor_n_5279: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4845,
        in1(1) => S4832,
        out1 => S4846
    );
nand_n_5280: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4846,
        in1(1) => S4831,
        out1 => S4848
    );
nand_n_5281: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4796,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S4849
    );
nand_n_5282: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4795,
        in1(1) => S5926,
        out1 => S4850
    );
notg_5283: ENTITY WORK.notg
    PORT MAP (
        in1 => S4850,
        out1 => S4851
    );
nand_n_5284: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4849,
        in1(1) => S4637,
        out1 => S4852
    );
nor_n_5285: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4852,
        in1(1) => S4851,
        out1 => S4853
    );
nor_n_5286: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4853,
        in1(1) => S4822,
        out1 => S4854
    );
nor_n_5287: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4848,
        in1(1) => S4829,
        out1 => S4855
    );
nand_n_5288: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4855,
        in1(1) => S4854,
        out1 => new_datapath_indatatrf_5
    );
nand_n_5289: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4533,
        in1(1) => S4482,
        out1 => S4856
    );
nand_n_5290: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4856,
        in1(1) => S4623,
        out1 => S4858
    );
nor_n_5291: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4858,
        in1(1) => S4534,
        out1 => S4859
    );
nor_n_5292: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4830,
        in1(1) => S4826,
        out1 => S4860
    );
nand_n_5293: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4860,
        in1(1) => S4483,
        out1 => S4861
    );
nor_n_5294: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4860,
        in1(1) => S4483,
        out1 => S4862
    );
notg_5295: ENTITY WORK.notg
    PORT MAP (
        in1 => S4862,
        out1 => S4863
    );
nor_n_5296: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4862,
        in1(1) => S4626,
        out1 => S4864
    );
nand_n_5297: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4864,
        in1(1) => S4861,
        out1 => S4865
    );
nand_n_5298: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4850,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S4866
    );
nor_n_5299: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4850,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S4867
    );
nor_n_5300: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4867,
        in1(1) => S4638,
        out1 => S4869
    );
nand_n_5301: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4869,
        in1(1) => S4866,
        out1 => S4870
    );
nor_n_5302: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4630,
        in1(1) => S4480,
        out1 => S4871
    );
nand_n_5303: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4633,
        in1(1) => S4472,
        out1 => S4872
    );
nor_n_5304: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4661,
        in1(1) => S3511,
        out1 => S4873
    );
nand_n_5305: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4648,
        in1(1) => new_datapath_shiftunit_2373_A,
        out1 => S4874
    );
nor_n_5306: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4670,
        in1(1) => S6179,
        out1 => S4875
    );
nand_n_5307: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => new_datapath_multdivunit_outmdu1_6,
        out1 => S4876
    );
nand_n_5308: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6215,
        in1(1) => new_datapath_databusin_6,
        out1 => S4877
    );
nand_n_5309: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4144,
        in1(1) => new_datapath_multdivunit_outmdu2_6,
        out1 => S4878
    );
nand_n_5310: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4878,
        in1(1) => S4877,
        out1 => S4880
    );
notg_5311: ENTITY WORK.notg
    PORT MAP (
        in1 => S4880,
        out1 => S4881
    );
nand_n_5312: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4881,
        in1(1) => S4876,
        out1 => S4882
    );
nor_n_5313: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4882,
        in1(1) => S4875,
        out1 => S4883
    );
nand_n_5314: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4883,
        in1(1) => S4874,
        out1 => S4884
    );
nor_n_5315: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4884,
        in1(1) => S4873,
        out1 => S4885
    );
nand_n_5316: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4885,
        in1(1) => S4872,
        out1 => S4886
    );
nor_n_5317: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4886,
        in1(1) => S4871,
        out1 => S4887
    );
nand_n_5318: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4887,
        in1(1) => S4870,
        out1 => S4888
    );
nor_n_5319: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4888,
        in1(1) => S4859,
        out1 => S4889
    );
nand_n_5320: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4889,
        in1(1) => S4865,
        out1 => new_datapath_indatatrf_6
    );
nor_n_5321: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4535,
        in1(1) => S4321,
        out1 => S4891
    );
nor_n_5322: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4536,
        in1(1) => S4320,
        out1 => S4892
    );
nor_n_5323: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4892,
        in1(1) => S4891,
        out1 => S4893
    );
nor_n_5324: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4893,
        in1(1) => S4624,
        out1 => S4894
    );
nand_n_5325: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4863,
        in1(1) => S4480,
        out1 => S4895
    );
nor_n_5326: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4895,
        in1(1) => S4320,
        out1 => S4896
    );
nand_n_5327: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4895,
        in1(1) => S4320,
        out1 => S4897
    );
notg_5328: ENTITY WORK.notg
    PORT MAP (
        in1 => S4897,
        out1 => S4898
    );
nor_n_5329: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4898,
        in1(1) => S4896,
        out1 => S4899
    );
nand_n_5330: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4899,
        in1(1) => S4625,
        out1 => S4901
    );
nor_n_5331: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4630,
        in1(1) => S4316,
        out1 => S4902
    );
nand_n_5332: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4633,
        in1(1) => S4309,
        out1 => S4903
    );
nor_n_5333: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4661,
        in1(1) => S3522,
        out1 => S4904
    );
nand_n_5334: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4648,
        in1(1) => new_datapath_shiftunit_2391_A,
        out1 => S4905
    );
notg_5335: ENTITY WORK.notg
    PORT MAP (
        in1 => S4905,
        out1 => S4906
    );
nor_n_5336: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4670,
        in1(1) => S6193,
        out1 => S4907
    );
nand_n_5337: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => new_datapath_multdivunit_outmdu1_7,
        out1 => S4908
    );
nand_n_5338: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6215,
        in1(1) => new_datapath_databusin_7,
        out1 => S4909
    );
nand_n_5339: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4144,
        in1(1) => new_datapath_multdivunit_outmdu2_7,
        out1 => S4910
    );
nand_n_5340: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4910,
        in1(1) => S4908,
        out1 => S4912
    );
nor_n_5341: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4912,
        in1(1) => S4907,
        out1 => S4913
    );
nand_n_5342: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4913,
        in1(1) => S4909,
        out1 => S4914
    );
nor_n_5343: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4914,
        in1(1) => S4906,
        out1 => S4915
    );
nor_n_5344: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4867,
        in1(1) => S5907,
        out1 => S4916
    );
nand_n_5345: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4867,
        in1(1) => S5907,
        out1 => S4917
    );
nand_n_5346: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4917,
        in1(1) => S4637,
        out1 => S4918
    );
nor_n_5347: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4918,
        in1(1) => S4916,
        out1 => S4919
    );
nand_n_5348: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4915,
        in1(1) => S4903,
        out1 => S4920
    );
nor_n_5349: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4920,
        in1(1) => S4902,
        out1 => S4921
    );
nor_n_5350: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4919,
        in1(1) => S4904,
        out1 => S4923
    );
nand_n_5351: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4923,
        in1(1) => S4921,
        out1 => S4924
    );
nor_n_5352: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4924,
        in1(1) => S4894,
        out1 => S4925
    );
nand_n_5353: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4925,
        in1(1) => S4901,
        out1 => new_datapath_indatatrf_7
    );
nand_n_5354: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4538,
        in1(1) => S4447,
        out1 => S4926
    );
nand_n_5355: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4926,
        in1(1) => S4623,
        out1 => S4927
    );
nor_n_5356: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4927,
        in1(1) => S4539,
        out1 => S4928
    );
nor_n_5357: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4895,
        in1(1) => S4315,
        out1 => S4929
    );
nor_n_5358: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4929,
        in1(1) => S4317,
        out1 => S4930
    );
nand_n_5359: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4930,
        in1(1) => S4447,
        out1 => S4931
    );
nor_n_5360: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4930,
        in1(1) => S4447,
        out1 => S4933
    );
nor_n_5361: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4933,
        in1(1) => S4626,
        out1 => S4934
    );
nand_n_5362: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4934,
        in1(1) => S4931,
        out1 => S4935
    );
nand_n_5363: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4917,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S4936
    );
nor_n_5364: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4917,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S4937
    );
nor_n_5365: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4937,
        in1(1) => S4638,
        out1 => S4938
    );
nand_n_5366: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4938,
        in1(1) => S4936,
        out1 => S4939
    );
nor_n_5367: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4661,
        in1(1) => S3533,
        out1 => S4940
    );
nand_n_5368: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4648,
        in1(1) => new_datapath_shiftunit_2409_A,
        out1 => S4941
    );
nand_n_5369: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4629,
        in1(1) => S4444,
        out1 => S4942
    );
nand_n_5370: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4633,
        in1(1) => S4389,
        out1 => S4944
    );
nor_n_5371: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4670,
        in1(1) => S6205,
        out1 => S4945
    );
nand_n_5372: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => new_datapath_multdivunit_outmdu1_8,
        out1 => S4946
    );
nand_n_5373: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6215,
        in1(1) => new_datapath_databusin_8,
        out1 => S4947
    );
nand_n_5374: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4144,
        in1(1) => new_datapath_multdivunit_outmdu2_8,
        out1 => S4948
    );
nand_n_5375: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4947,
        in1(1) => S4944,
        out1 => S4949
    );
nand_n_5376: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4948,
        in1(1) => S4946,
        out1 => S4950
    );
nor_n_5377: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4950,
        in1(1) => S4945,
        out1 => S4951
    );
nand_n_5378: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4951,
        in1(1) => S4942,
        out1 => S4952
    );
nor_n_5379: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4952,
        in1(1) => S4949,
        out1 => S4953
    );
nand_n_5380: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4953,
        in1(1) => S4941,
        out1 => S4955
    );
nor_n_5381: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4955,
        in1(1) => S4940,
        out1 => S4956
    );
nand_n_5382: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4956,
        in1(1) => S4939,
        out1 => S4957
    );
nor_n_5383: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4957,
        in1(1) => S4928,
        out1 => S4958
    );
nand_n_5384: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4958,
        in1(1) => S4935,
        out1 => new_datapath_indatatrf_8
    );
nor_n_5385: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4542,
        in1(1) => S4455,
        out1 => S4959
    );
nor_n_5386: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4543,
        in1(1) => S4456,
        out1 => S4960
    );
nor_n_5387: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4960,
        in1(1) => S4959,
        out1 => S4961
    );
nand_n_5388: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4961,
        in1(1) => S4623,
        out1 => S4962
    );
nand_n_5389: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4931,
        in1(1) => S4442,
        out1 => S4963
    );
nor_n_5390: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4963,
        in1(1) => S4456,
        out1 => S4965
    );
nand_n_5391: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4963,
        in1(1) => S4456,
        out1 => S4966
    );
nand_n_5392: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4966,
        in1(1) => S4625,
        out1 => S4967
    );
nor_n_5393: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4967,
        in1(1) => S4965,
        out1 => S4968
    );
nor_n_5394: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4937,
        in1(1) => S3336,
        out1 => S4969
    );
nand_n_5395: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4937,
        in1(1) => S3336,
        out1 => S4970
    );
nand_n_5396: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4970,
        in1(1) => S4637,
        out1 => S4971
    );
nor_n_5397: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4971,
        in1(1) => S4969,
        out1 => S4972
    );
nor_n_5398: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4661,
        in1(1) => S3544,
        out1 => S4973
    );
nand_n_5399: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4648,
        in1(1) => new_datapath_shiftunit_2427_A,
        out1 => S4974
    );
nand_n_5400: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4450,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S4976
    );
nor_n_5401: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4976,
        in1(1) => S4630,
        out1 => S4977
    );
nor_n_5402: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4285,
        in1(1) => new_controller_fib_1,
        out1 => S4978
    );
nor_n_5403: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4978,
        in1(1) => S4384,
        out1 => S4979
    );
nor_n_5404: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4979,
        in1(1) => S4306,
        out1 => S4980
    );
nor_n_5405: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4980,
        in1(1) => S4634,
        out1 => S4981
    );
nand_n_5406: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4669,
        in1(1) => S93,
        out1 => S4982
    );
nand_n_5407: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => new_datapath_multdivunit_outmdu1_9,
        out1 => S4983
    );
nand_n_5408: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6215,
        in1(1) => new_datapath_databusin_9,
        out1 => S4984
    );
nand_n_5409: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4144,
        in1(1) => new_datapath_multdivunit_outmdu2_9,
        out1 => S4985
    );
nand_n_5410: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4985,
        in1(1) => S4983,
        out1 => S4987
    );
nor_n_5411: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4987,
        in1(1) => S4981,
        out1 => S4988
    );
nand_n_5412: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4988,
        in1(1) => S4982,
        out1 => S4989
    );
nor_n_5413: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4989,
        in1(1) => S4977,
        out1 => S4990
    );
nand_n_5414: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4990,
        in1(1) => S4984,
        out1 => S4991
    );
nor_n_5415: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4991,
        in1(1) => S4973,
        out1 => S4992
    );
nand_n_5416: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4992,
        in1(1) => S4974,
        out1 => S4993
    );
nor_n_5417: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4993,
        in1(1) => S4972,
        out1 => S4994
    );
notg_5418: ENTITY WORK.notg
    PORT MAP (
        in1 => S4994,
        out1 => S4995
    );
nor_n_5419: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4995,
        in1(1) => S4968,
        out1 => S4996
    );
nand_n_5420: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4996,
        in1(1) => S4962,
        out1 => new_datapath_indatatrf_9
    );
nand_n_5421: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4545,
        in1(1) => S4438,
        out1 => S4998
    );
nor_n_5422: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4624,
        in1(1) => S4546,
        out1 => S4999
    );
nand_n_5423: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4999,
        in1(1) => S4998,
        out1 => S5000
    );
nand_n_5424: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4976,
        in1(1) => S4966,
        out1 => S5001
    );
nor_n_5425: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5001,
        in1(1) => S4438,
        out1 => S5002
    );
nand_n_5426: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5001,
        in1(1) => S4438,
        out1 => S5003
    );
nand_n_5427: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5003,
        in1(1) => S4625,
        out1 => S5004
    );
nor_n_5428: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5004,
        in1(1) => S5002,
        out1 => S5005
    );
nand_n_5429: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4970,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S5006
    );
nor_n_5430: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4970,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S5008
    );
notg_5431: ENTITY WORK.notg
    PORT MAP (
        in1 => S5008,
        out1 => S5009
    );
nor_n_5432: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5008,
        in1(1) => S4638,
        out1 => S5010
    );
nand_n_5433: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5010,
        in1(1) => S5006,
        out1 => S5011
    );
nor_n_5434: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4661,
        in1(1) => S3554,
        out1 => S5012
    );
nand_n_5435: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4648,
        in1(1) => new_datapath_shiftunit_2445_A,
        out1 => S5013
    );
nor_n_5436: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4630,
        in1(1) => S4435,
        out1 => S5014
    );
nand_n_5437: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4669,
        in1(1) => S107,
        out1 => S5015
    );
nor_n_5438: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4285,
        in1(1) => new_controller_fib_2,
        out1 => S5016
    );
nor_n_5439: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5016,
        in1(1) => S4384,
        out1 => S5017
    );
nor_n_5440: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5017,
        in1(1) => S4306,
        out1 => S5019
    );
nor_n_5441: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5019,
        in1(1) => S4634,
        out1 => S5020
    );
nand_n_5442: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4144,
        in1(1) => new_datapath_multdivunit_outmdu2_10,
        out1 => S5021
    );
nand_n_5443: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => new_datapath_multdivunit_outmdu1_10,
        out1 => S5022
    );
nand_n_5444: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6215,
        in1(1) => new_datapath_databusin_10,
        out1 => S5023
    );
nand_n_5445: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5023,
        in1(1) => S5022,
        out1 => S5024
    );
notg_5446: ENTITY WORK.notg
    PORT MAP (
        in1 => S5024,
        out1 => S5025
    );
nand_n_5447: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5025,
        in1(1) => S5021,
        out1 => S5026
    );
nor_n_5448: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5026,
        in1(1) => S5020,
        out1 => S5027
    );
nand_n_5449: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5027,
        in1(1) => S5015,
        out1 => S5028
    );
nor_n_5450: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5028,
        in1(1) => S5014,
        out1 => S5030
    );
nand_n_5451: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5030,
        in1(1) => S5013,
        out1 => S5031
    );
nor_n_5452: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5031,
        in1(1) => S5012,
        out1 => S5032
    );
nand_n_5453: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5032,
        in1(1) => S5011,
        out1 => S5033
    );
nor_n_5454: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5033,
        in1(1) => S5005,
        out1 => S5034
    );
nand_n_5455: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5034,
        in1(1) => S5000,
        out1 => new_datapath_indatatrf_10
    );
nand_n_5456: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4547,
        in1(1) => S4467,
        out1 => S5035
    );
nor_n_5457: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4547,
        in1(1) => S4467,
        out1 => S5036
    );
notg_5458: ENTITY WORK.notg
    PORT MAP (
        in1 => S5036,
        out1 => S5037
    );
nand_n_5459: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5037,
        in1(1) => S5035,
        out1 => S5038
    );
nor_n_5460: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5038,
        in1(1) => S4624,
        out1 => S5040
    );
nand_n_5461: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5003,
        in1(1) => S4435,
        out1 => S5041
    );
nor_n_5462: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5041,
        in1(1) => S4467,
        out1 => S5042
    );
notg_5463: ENTITY WORK.notg
    PORT MAP (
        in1 => S5042,
        out1 => S5043
    );
nand_n_5464: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5041,
        in1(1) => S4467,
        out1 => S5044
    );
nand_n_5465: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5044,
        in1(1) => S5043,
        out1 => S5045
    );
nor_n_5466: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5045,
        in1(1) => S4626,
        out1 => S5046
    );
nor_n_5467: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4661,
        in1(1) => S3565,
        out1 => S5047
    );
nand_n_5468: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4648,
        in1(1) => new_datapath_shiftunit_2463_A,
        out1 => S5048
    );
nand_n_5469: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4629,
        in1(1) => S4464,
        out1 => S5049
    );
nor_n_5470: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4670,
        in1(1) => S122,
        out1 => S5051
    );
nor_n_5471: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4285,
        in1(1) => new_controller_fib_3,
        out1 => S5052
    );
nor_n_5472: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5052,
        in1(1) => S4384,
        out1 => S5053
    );
nor_n_5473: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5053,
        in1(1) => S4306,
        out1 => S5054
    );
nor_n_5474: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5054,
        in1(1) => S4634,
        out1 => S5055
    );
nand_n_5475: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4144,
        in1(1) => new_datapath_multdivunit_outmdu2_11,
        out1 => S5056
    );
nand_n_5476: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6215,
        in1(1) => new_datapath_databusin_11,
        out1 => S5057
    );
nand_n_5477: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5057,
        in1(1) => S5056,
        out1 => S5058
    );
nand_n_5478: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => new_datapath_multdivunit_outmdu1_11,
        out1 => S5059
    );
nor_n_5479: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5055,
        in1(1) => S5051,
        out1 => S5060
    );
nand_n_5480: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5059,
        in1(1) => S5049,
        out1 => S5062
    );
nor_n_5481: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5062,
        in1(1) => S5058,
        out1 => S5063
    );
nand_n_5482: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5063,
        in1(1) => S5048,
        out1 => S5064
    );
nor_n_5483: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5064,
        in1(1) => S5047,
        out1 => S5065
    );
nand_n_5484: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5065,
        in1(1) => S5060,
        out1 => S5066
    );
nand_n_5485: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5009,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S5067
    );
nand_n_5486: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5008,
        in1(1) => S3357,
        out1 => S5068
    );
nand_n_5487: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5068,
        in1(1) => S5067,
        out1 => S5069
    );
nor_n_5488: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5069,
        in1(1) => S4638,
        out1 => S5070
    );
nor_n_5489: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5066,
        in1(1) => S5040,
        out1 => S5071
    );
nor_n_5490: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5070,
        in1(1) => S5046,
        out1 => S5073
    );
nand_n_5491: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5073,
        in1(1) => S5071,
        out1 => new_datapath_indatatrf_11
    );
nand_n_5492: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4549,
        in1(1) => S4427,
        out1 => S5074
    );
nor_n_5493: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4549,
        in1(1) => S4427,
        out1 => S5075
    );
notg_5494: ENTITY WORK.notg
    PORT MAP (
        in1 => S5075,
        out1 => S5076
    );
nor_n_5495: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5075,
        in1(1) => S4624,
        out1 => S5077
    );
nand_n_5496: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5077,
        in1(1) => S5074,
        out1 => S5078
    );
nor_n_5497: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5041,
        in1(1) => S4464,
        out1 => S5079
    );
nor_n_5498: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5079,
        in1(1) => S4466,
        out1 => S5080
    );
nor_n_5499: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5080,
        in1(1) => S4427,
        out1 => S5081
    );
nand_n_5500: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5080,
        in1(1) => S4427,
        out1 => S5083
    );
notg_5501: ENTITY WORK.notg
    PORT MAP (
        in1 => S5083,
        out1 => S5084
    );
nand_n_5502: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5083,
        in1(1) => S4625,
        out1 => S5085
    );
nor_n_5503: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5085,
        in1(1) => S5081,
        out1 => S5086
    );
nand_n_5504: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5068,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S5087
    );
nor_n_5505: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5068,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S5088
    );
notg_5506: ENTITY WORK.notg
    PORT MAP (
        in1 => S5088,
        out1 => S5089
    );
nor_n_5507: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5088,
        in1(1) => S4638,
        out1 => S5090
    );
nand_n_5508: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5090,
        in1(1) => S5087,
        out1 => S5091
    );
nor_n_5509: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4661,
        in1(1) => S3576,
        out1 => S5092
    );
nand_n_5510: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4648,
        in1(1) => new_datapath_shiftunit_2481_A,
        out1 => S5094
    );
nor_n_5511: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4670,
        in1(1) => S134,
        out1 => S5095
    );
nand_n_5512: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4629,
        in1(1) => S4424,
        out1 => S5096
    );
nor_n_5513: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4285,
        in1(1) => new_controller_fib_4,
        out1 => S5097
    );
nor_n_5514: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5097,
        in1(1) => S4384,
        out1 => S5098
    );
nor_n_5515: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5098,
        in1(1) => S4306,
        out1 => S5099
    );
nor_n_5516: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5099,
        in1(1) => S4634,
        out1 => S5100
    );
nand_n_5517: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4144,
        in1(1) => new_datapath_multdivunit_outmdu2_12,
        out1 => S5101
    );
nand_n_5518: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6215,
        in1(1) => new_datapath_databusin_12,
        out1 => S5102
    );
nand_n_5519: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => new_datapath_multdivunit_outmdu1_12,
        out1 => S5103
    );
nand_n_5520: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5103,
        in1(1) => S5102,
        out1 => S5105
    );
notg_5521: ENTITY WORK.notg
    PORT MAP (
        in1 => S5105,
        out1 => S5106
    );
nand_n_5522: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5106,
        in1(1) => S5101,
        out1 => S5107
    );
nor_n_5523: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5107,
        in1(1) => S5100,
        out1 => S5108
    );
nand_n_5524: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5108,
        in1(1) => S5096,
        out1 => S5109
    );
nor_n_5525: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5109,
        in1(1) => S5095,
        out1 => S5110
    );
nand_n_5526: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5110,
        in1(1) => S5094,
        out1 => S5111
    );
nor_n_5527: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5111,
        in1(1) => S5092,
        out1 => S5112
    );
nand_n_5528: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5112,
        in1(1) => S5091,
        out1 => S5113
    );
nor_n_5529: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5113,
        in1(1) => S5086,
        out1 => S5114
    );
nand_n_5530: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5114,
        in1(1) => S5078,
        out1 => new_datapath_indatatrf_12
    );
nand_n_5531: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5076,
        in1(1) => S4426,
        out1 => S5116
    );
nand_n_5532: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5116,
        in1(1) => S4418,
        out1 => S5117
    );
nor_n_5533: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5116,
        in1(1) => S4418,
        out1 => S5118
    );
nor_n_5534: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5118,
        in1(1) => S4624,
        out1 => S5119
    );
nand_n_5535: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5119,
        in1(1) => S5117,
        out1 => S5120
    );
nor_n_5536: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5084,
        in1(1) => S4424,
        out1 => S5121
    );
nor_n_5537: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5121,
        in1(1) => S4417,
        out1 => S5122
    );
nand_n_5538: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5121,
        in1(1) => S4417,
        out1 => S5123
    );
notg_5539: ENTITY WORK.notg
    PORT MAP (
        in1 => S5123,
        out1 => S5124
    );
nor_n_5540: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5124,
        in1(1) => S5122,
        out1 => S5126
    );
nor_n_5541: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5126,
        in1(1) => S4626,
        out1 => S5127
    );
nor_n_5542: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5088,
        in1(1) => S3379,
        out1 => S5128
    );
nor_n_5543: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5089,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S5129
    );
notg_5544: ENTITY WORK.notg
    PORT MAP (
        in1 => S5129,
        out1 => S5130
    );
nor_n_5545: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5129,
        in1(1) => S5128,
        out1 => S5131
    );
nand_n_5546: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5131,
        in1(1) => S4637,
        out1 => S5132
    );
nand_n_5547: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4660,
        in1(1) => new_datapath_shiftunit_2195_A,
        out1 => S5133
    );
nand_n_5548: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4648,
        in1(1) => new_datapath_shiftunit_2499_A,
        out1 => S5134
    );
nor_n_5549: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4670,
        in1(1) => S148,
        out1 => S5135
    );
nand_n_5550: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4629,
        in1(1) => S4416,
        out1 => S5137
    );
nor_n_5551: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4285,
        in1(1) => new_controller_234_B_0,
        out1 => S5138
    );
nor_n_5552: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5138,
        in1(1) => S4384,
        out1 => S5139
    );
nor_n_5553: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5139,
        in1(1) => S4306,
        out1 => S5140
    );
nor_n_5554: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5140,
        in1(1) => S4634,
        out1 => S5141
    );
nand_n_5555: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4144,
        in1(1) => new_datapath_multdivunit_outmdu2_13,
        out1 => S5142
    );
nand_n_5556: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => new_datapath_multdivunit_outmdu1_13,
        out1 => S5143
    );
nand_n_5557: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6215,
        in1(1) => new_datapath_databusin_13,
        out1 => S5144
    );
nand_n_5558: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5144,
        in1(1) => S5134,
        out1 => S5145
    );
nand_n_5559: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5143,
        in1(1) => S5142,
        out1 => S5146
    );
nor_n_5560: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5146,
        in1(1) => S5141,
        out1 => S5148
    );
nand_n_5561: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5148,
        in1(1) => S5137,
        out1 => S5149
    );
nor_n_5562: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5149,
        in1(1) => S5135,
        out1 => S5150
    );
nand_n_5563: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5150,
        in1(1) => S5133,
        out1 => S5151
    );
nor_n_5564: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5151,
        in1(1) => S5145,
        out1 => S5152
    );
nand_n_5565: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5152,
        in1(1) => S5132,
        out1 => S5153
    );
nor_n_5566: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5153,
        in1(1) => S5127,
        out1 => S5154
    );
nand_n_5567: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5154,
        in1(1) => S5120,
        out1 => new_datapath_indatatrf_13
    );
nand_n_5568: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5117,
        in1(1) => S4554,
        out1 => S5155
    );
nor_n_5569: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5155,
        in1(1) => S4409,
        out1 => S5156
    );
nand_n_5570: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5155,
        in1(1) => S4409,
        out1 => S5158
    );
nand_n_5571: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5158,
        in1(1) => S4623,
        out1 => S5159
    );
nor_n_5572: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5159,
        in1(1) => S5156,
        out1 => S5160
    );
nor_n_5573: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5121,
        in1(1) => S4415,
        out1 => S5161
    );
nor_n_5574: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5161,
        in1(1) => S4416,
        out1 => S5162
    );
nand_n_5575: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5162,
        in1(1) => S4409,
        out1 => S5163
    );
nor_n_5576: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5162,
        in1(1) => S4409,
        out1 => S5164
    );
nor_n_5577: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5164,
        in1(1) => S4626,
        out1 => S5165
    );
nand_n_5578: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5165,
        in1(1) => S5163,
        out1 => S5166
    );
nor_n_5579: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5130,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S5167
    );
nor_n_5580: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5129,
        in1(1) => S3390,
        out1 => S5169
    );
nor_n_5581: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5169,
        in1(1) => S5167,
        out1 => S5170
    );
nand_n_5582: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5170,
        in1(1) => S4637,
        out1 => S5171
    );
nand_n_5583: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4660,
        in1(1) => new_datapath_shiftunit_2213_A,
        out1 => S5172
    );
nand_n_5584: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4648,
        in1(1) => new_datapath_shiftunit_2517_A,
        out1 => S5173
    );
nand_n_5585: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4629,
        in1(1) => S4408,
        out1 => S5174
    );
nor_n_5586: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4285,
        in1(1) => new_controller_opcode_2,
        out1 => S5175
    );
nor_n_5587: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5175,
        in1(1) => S4384,
        out1 => S5176
    );
nor_n_5588: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5176,
        in1(1) => S4306,
        out1 => S5177
    );
nor_n_5589: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5177,
        in1(1) => S4634,
        out1 => S5178
    );
nand_n_5590: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => new_datapath_multdivunit_outmdu1_14,
        out1 => S5180
    );
nor_n_5591: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3740,
        in1(1) => S3106,
        out1 => S5181
    );
nand_n_5592: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4144,
        in1(1) => new_datapath_multdivunit_outmdu2_14,
        out1 => S5182
    );
nand_n_5593: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5182,
        in1(1) => S5180,
        out1 => S5183
    );
nor_n_5594: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5183,
        in1(1) => S5178,
        out1 => S5184
    );
nand_n_5595: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5184,
        in1(1) => S5174,
        out1 => S5185
    );
nor_n_5596: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5185,
        in1(1) => S5181,
        out1 => S5186
    );
nand_n_5597: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5186,
        in1(1) => S5173,
        out1 => S5187
    );
nand_n_5598: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4669,
        in1(1) => S161,
        out1 => S5188
    );
nand_n_5599: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5188,
        in1(1) => S5172,
        out1 => S5189
    );
nor_n_5600: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5189,
        in1(1) => S5187,
        out1 => S5191
    );
nand_n_5601: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5191,
        in1(1) => S5171,
        out1 => S5192
    );
nor_n_5602: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5192,
        in1(1) => S5160,
        out1 => S5193
    );
nand_n_5603: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5193,
        in1(1) => S5166,
        out1 => new_datapath_indatatrf_14
    );
nand_n_5604: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5158,
        in1(1) => S4406,
        out1 => S5194
    );
nand_n_5605: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5194,
        in1(1) => S4401,
        out1 => S5195
    );
nor_n_5606: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5194,
        in1(1) => S4401,
        out1 => S5196
    );
nor_n_5607: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5196,
        in1(1) => S4624,
        out1 => S5197
    );
nand_n_5608: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5197,
        in1(1) => S5195,
        out1 => S5198
    );
nor_n_5609: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5164,
        in1(1) => S4408,
        out1 => S5199
    );
nand_n_5610: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5199,
        in1(1) => S4401,
        out1 => S5201
    );
nor_n_5611: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5199,
        in1(1) => S4401,
        out1 => S5202
    );
nand_n_5612: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5201,
        in1(1) => S4625,
        out1 => S5203
    );
nor_n_5613: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5203,
        in1(1) => S5202,
        out1 => S5204
    );
nor_n_5614: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4670,
        in1(1) => S6075,
        out1 => S5205
    );
nand_n_5615: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4660,
        in1(1) => new_datapath_shiftunit_2231_A,
        out1 => S5206
    );
nand_n_5616: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4648,
        in1(1) => new_datapath_shiftunit_2534_A,
        out1 => S5207
    );
nand_n_5617: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4629,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S5208
    );
nor_n_5618: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5208,
        in1(1) => S4394,
        out1 => S5209
    );
nor_n_5619: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4383,
        in1(1) => S4306,
        out1 => S5210
    );
nor_n_5620: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5210,
        in1(1) => S4634,
        out1 => S5212
    );
nor_n_5621: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4155,
        in1(1) => S2581,
        out1 => S5213
    );
nor_n_5622: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S3740,
        in1(1) => S2603,
        out1 => S5214
    );
nand_n_5623: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => new_datapath_multdivunit_outmdu1_15,
        out1 => S5215
    );
nor_n_5624: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5213,
        in1(1) => S5212,
        out1 => S5216
    );
nand_n_5625: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5216,
        in1(1) => S5206,
        out1 => S5217
    );
nor_n_5626: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5214,
        in1(1) => S5205,
        out1 => S5218
    );
nand_n_5627: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5215,
        in1(1) => S5207,
        out1 => S5219
    );
nor_n_5628: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5219,
        in1(1) => S5209,
        out1 => S5220
    );
nand_n_5629: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5220,
        in1(1) => S5218,
        out1 => S5221
    );
nor_n_5630: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5221,
        in1(1) => S5217,
        out1 => S5223
    );
nand_n_5631: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5167,
        in1(1) => S3401,
        out1 => S5224
    );
nor_n_5632: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5167,
        in1(1) => S3401,
        out1 => S5225
    );
nor_n_5633: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5225,
        in1(1) => S4638,
        out1 => S5226
    );
nand_n_5634: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5226,
        in1(1) => S5224,
        out1 => S5227
    );
nand_n_5635: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5227,
        in1(1) => S5223,
        out1 => S5228
    );
nor_n_5636: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5228,
        in1(1) => S5204,
        out1 => S5229
    );
nand_n_5637: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5229,
        in1(1) => S5198,
        out1 => new_datapath_indatatrf_15
    );
nand_n_5638: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_muxmem_in2_0,
        out1 => S5230
    );
nand_n_5639: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3708,
        in1(1) => new_datapath_adr_outreg_0,
        out1 => S5231
    );
nand_n_5640: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5231,
        in1(1) => S5230,
        out1 => new_datapath_addrbus_0
    );
nand_n_5641: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_muxmem_in2_1,
        out1 => S5233
    );
nand_n_5642: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3708,
        in1(1) => new_datapath_adr_outreg_1,
        out1 => S5234
    );
nand_n_5643: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5234,
        in1(1) => S5233,
        out1 => new_datapath_addrbus_1
    );
nand_n_5644: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_muxmem_in2_2,
        out1 => S5235
    );
nand_n_5645: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3708,
        in1(1) => new_datapath_adr_outreg_2,
        out1 => S5236
    );
nand_n_5646: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5236,
        in1(1) => S5235,
        out1 => new_datapath_addrbus_2
    );
nand_n_5647: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_muxmem_in2_3,
        out1 => S5237
    );
nand_n_5648: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3708,
        in1(1) => new_datapath_adr_outreg_3,
        out1 => S5238
    );
nand_n_5649: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5238,
        in1(1) => S5237,
        out1 => new_datapath_addrbus_3
    );
nand_n_5650: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_muxmem_in2_4,
        out1 => S5240
    );
nand_n_5651: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3708,
        in1(1) => new_datapath_adr_outreg_4,
        out1 => S5241
    );
nand_n_5652: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5241,
        in1(1) => S5240,
        out1 => new_datapath_addrbus_4
    );
nand_n_5653: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_muxmem_in2_5,
        out1 => S5242
    );
nand_n_5654: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3708,
        in1(1) => new_datapath_adr_outreg_5,
        out1 => S5243
    );
nand_n_5655: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5243,
        in1(1) => S5242,
        out1 => new_datapath_addrbus_5
    );
nand_n_5656: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_muxmem_in2_6,
        out1 => S5244
    );
nand_n_5657: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3708,
        in1(1) => new_datapath_adr_outreg_6,
        out1 => S5245
    );
nand_n_5658: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5245,
        in1(1) => S5244,
        out1 => new_datapath_addrbus_6
    );
nand_n_5659: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_muxmem_in2_7,
        out1 => S5246
    );
nand_n_5660: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3708,
        in1(1) => new_datapath_adr_outreg_7,
        out1 => S5248
    );
nand_n_5661: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5248,
        in1(1) => S5246,
        out1 => new_datapath_addrbus_7
    );
nand_n_5662: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_muxmem_in2_8,
        out1 => S5249
    );
nand_n_5663: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3708,
        in1(1) => new_datapath_adr_outreg_8,
        out1 => S5250
    );
nand_n_5664: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5250,
        in1(1) => S5249,
        out1 => new_datapath_addrbus_8
    );
nand_n_5665: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_muxmem_in2_9,
        out1 => S5251
    );
nand_n_5666: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3708,
        in1(1) => new_datapath_adr_outreg_9,
        out1 => S5252
    );
nand_n_5667: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5252,
        in1(1) => S5251,
        out1 => new_datapath_addrbus_9
    );
nand_n_5668: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_muxmem_in2_10,
        out1 => S5253
    );
nand_n_5669: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3708,
        in1(1) => new_datapath_adr_outreg_10,
        out1 => S5254
    );
nand_n_5670: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5254,
        in1(1) => S5253,
        out1 => new_datapath_addrbus_10
    );
nand_n_5671: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_muxmem_in2_11,
        out1 => S5256
    );
nand_n_5672: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3708,
        in1(1) => new_datapath_adr_outreg_11,
        out1 => S5257
    );
nand_n_5673: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5257,
        in1(1) => S5256,
        out1 => new_datapath_addrbus_11
    );
nand_n_5674: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_muxmem_in2_12,
        out1 => S5258
    );
nand_n_5675: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3708,
        in1(1) => new_datapath_adr_outreg_12,
        out1 => S5259
    );
nand_n_5676: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5259,
        in1(1) => S5258,
        out1 => new_datapath_addrbus_12
    );
nand_n_5677: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_muxmem_in2_13,
        out1 => S5260
    );
nand_n_5678: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3708,
        in1(1) => new_datapath_adr_outreg_13,
        out1 => S5261
    );
nand_n_5679: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5261,
        in1(1) => S5260,
        out1 => new_datapath_addrbus_13
    );
nand_n_5680: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_muxmem_in2_14,
        out1 => S5263
    );
nand_n_5681: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3708,
        in1(1) => new_datapath_adr_outreg_14,
        out1 => S5264
    );
nand_n_5682: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5264,
        in1(1) => S5263,
        out1 => new_datapath_addrbus_14
    );
nand_n_5683: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_controller_1133_S_0,
        in1(1) => new_datapath_muxmem_in2_15,
        out1 => S5265
    );
nand_n_5684: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S3708,
        in1(1) => new_datapath_adr_outreg_15,
        out1 => S5266
    );
nand_n_5685: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5266,
        in1(1) => S5265,
        out1 => new_datapath_addrbus_15
    );
nor_n_5686: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S6086,
        in1(1) => S6215,
        out1 => S5267
    );
nand_n_5687: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5267,
        in1(1) => S4610,
        out1 => S5268
    );
notg_5688: ENTITY WORK.notg
    PORT MAP (
        in1 => S5268,
        out1 => S5269
    );
nand_n_5689: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5268,
        in1(1) => new_datapath_instruction_0,
        out1 => S5270
    );
nand_n_5690: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4144,
        in1(1) => S2964,
        out1 => S5272
    );
nand_n_5691: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5272,
        in1(1) => S5270,
        out1 => new_datapath_muxrd_outmux_0
    );
nor_n_5692: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => new_datapath_instruction_1,
        in1(1) => new_datapath_instruction_0,
        out1 => S5273
    );
nand_n_5693: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5268,
        in1(1) => new_datapath_instruction_1,
        out1 => S5274
    );
nand_n_5694: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => new_datapath_instruction_1,
        in1(1) => new_datapath_instruction_0,
        out1 => S5275
    );
notg_5695: ENTITY WORK.notg
    PORT MAP (
        in1 => S5275,
        out1 => S5276
    );
nor_n_5696: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5273,
        in1(1) => S4155,
        out1 => S5277
    );
nand_n_5697: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5277,
        in1(1) => S5275,
        out1 => S5278
    );
nand_n_5698: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5278,
        in1(1) => S5274,
        out1 => new_datapath_muxrd_outmux_1
    );
nand_n_5699: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5276,
        in1(1) => new_datapath_instruction_2,
        out1 => S5279
    );
nand_n_5700: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5279,
        in1(1) => S4144,
        out1 => S5281
    );
notg_5701: ENTITY WORK.notg
    PORT MAP (
        in1 => S5281,
        out1 => S5282
    );
nor_n_5702: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5282,
        in1(1) => S5268,
        out1 => S5283
    );
nand_n_5703: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5281,
        in1(1) => S5269,
        out1 => S5284
    );
nor_n_5704: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5281,
        in1(1) => S5275,
        out1 => S5285
    );
nor_n_5705: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5285,
        in1(1) => new_datapath_instruction_2,
        out1 => S5286
    );
nor_n_5706: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5286,
        in1(1) => S5283,
        out1 => new_datapath_muxrd_outmux_2
    );
nor_n_5707: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5279,
        in1(1) => S4155,
        out1 => S5287
    );
nor_n_5708: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5287,
        in1(1) => new_datapath_instruction_3,
        out1 => S5288
    );
nor_n_5709: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5284,
        in1(1) => S2975,
        out1 => S5289
    );
nor_n_5710: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5289,
        in1(1) => S5288,
        out1 => new_datapath_muxrd_outmux_3
    );
nor_n_5711: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S270,
        in1(1) => S5693,
        out1 => S5291
    );
nand_n_5712: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S271,
        in1(1) => S5683,
        out1 => S5292
    );
nor_n_5713: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5125,
        in1(1) => S2985,
        out1 => S5293
    );
nand_n_5714: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5115,
        in1(1) => new_controller_fib_0,
        out1 => S5294
    );
nor_n_5715: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5293,
        in1(1) => S5291,
        out1 => S5295
    );
nand_n_5716: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5294,
        in1(1) => S5292,
        out1 => S5296
    );
nor_n_5717: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S256,
        in1(1) => S5693,
        out1 => S5297
    );
nand_n_5718: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S257,
        in1(1) => S5683,
        out1 => S5298
    );
nor_n_5719: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5125,
        in1(1) => S3007,
        out1 => S5299
    );
nand_n_5720: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5115,
        in1(1) => new_controller_fib_2,
        out1 => S5301
    );
nor_n_5721: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5299,
        in1(1) => S5297,
        out1 => S5302
    );
nand_n_5722: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5301,
        in1(1) => S5298,
        out1 => S5303
    );
nor_n_5723: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S264,
        in1(1) => S5693,
        out1 => S5304
    );
nand_n_5724: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S265,
        in1(1) => S5683,
        out1 => S5305
    );
nor_n_5725: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5125,
        in1(1) => S2996,
        out1 => S5306
    );
nand_n_5726: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5115,
        in1(1) => new_controller_fib_1,
        out1 => S5307
    );
nor_n_5727: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5306,
        in1(1) => S5304,
        out1 => S5308
    );
nand_n_5728: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5307,
        in1(1) => S5305,
        out1 => S5309
    );
nor_n_5729: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S248,
        in1(1) => S5693,
        out1 => S5310
    );
nand_n_5730: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S249,
        in1(1) => S5683,
        out1 => S5312
    );
nor_n_5731: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5125,
        in1(1) => S3018,
        out1 => S5313
    );
nand_n_5732: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5115,
        in1(1) => new_controller_fib_3,
        out1 => S5314
    );
nor_n_5733: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5313,
        in1(1) => S5310,
        out1 => S5315
    );
nand_n_5734: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5314,
        in1(1) => S5312,
        out1 => S5316
    );
nor_n_5735: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5316,
        in1(1) => S5303,
        out1 => S5317
    );
nand_n_5736: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5315,
        in1(1) => S5302,
        out1 => S5318
    );
nor_n_5737: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5318,
        in1(1) => S5309,
        out1 => S5319
    );
nor_n_5738: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5309,
        in1(1) => S5296,
        out1 => S5320
    );
nand_n_5739: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5308,
        in1(1) => S5295,
        out1 => S5321
    );
nor_n_5740: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5321,
        in1(1) => S5318,
        out1 => S5323
    );
nand_n_5741: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5320,
        in1(1) => S5317,
        out1 => S5324
    );
nand_n_5742: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5323,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S5325
    );
notg_5743: ENTITY WORK.notg
    PORT MAP (
        in1 => S5325,
        out1 => new_datapath_shiftunit_2265_A
    );
nor_n_5744: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5315,
        in1(1) => S5303,
        out1 => S5326
    );
nand_n_5745: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5316,
        in1(1) => S5302,
        out1 => S5327
    );
nor_n_5746: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5327,
        in1(1) => S5321,
        out1 => S5328
    );
nand_n_5747: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5326,
        in1(1) => S5320,
        out1 => S5329
    );
nand_n_5748: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5328,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S5330
    );
nor_n_5749: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5308,
        in1(1) => S5295,
        out1 => S5331
    );
nand_n_5750: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5309,
        in1(1) => S5296,
        out1 => S5333
    );
nor_n_5751: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5316,
        in1(1) => S5302,
        out1 => S5334
    );
nand_n_5752: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5315,
        in1(1) => S5303,
        out1 => S5335
    );
nor_n_5753: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5335,
        in1(1) => S5333,
        out1 => S5336
    );
nand_n_5754: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5334,
        in1(1) => S5331,
        out1 => S5337
    );
nand_n_5755: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5336,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S5338
    );
nor_n_5756: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5309,
        in1(1) => S5295,
        out1 => S5339
    );
nand_n_5757: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5308,
        in1(1) => S5296,
        out1 => S5340
    );
nor_n_5758: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5315,
        in1(1) => S5302,
        out1 => S5341
    );
nand_n_5759: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5316,
        in1(1) => S5303,
        out1 => S5342
    );
nor_n_5760: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5342,
        in1(1) => S5340,
        out1 => S5344
    );
nand_n_5761: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5344,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S5345
    );
nor_n_5762: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5340,
        in1(1) => S5327,
        out1 => S5346
    );
nand_n_5763: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5346,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S5347
    );
nand_n_5764: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5347,
        in1(1) => S5345,
        out1 => S5348
    );
nor_n_5765: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5340,
        in1(1) => S5335,
        out1 => S5349
    );
nand_n_5766: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5349,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S5350
    );
nor_n_5767: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5342,
        in1(1) => S3401,
        out1 => S5351
    );
nand_n_5768: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5351,
        in1(1) => S5331,
        out1 => S5352
    );
nor_n_5769: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5333,
        in1(1) => S5327,
        out1 => S5353
    );
nand_n_5770: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5353,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S5355
    );
nor_n_5771: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5308,
        in1(1) => S5296,
        out1 => S5356
    );
nand_n_5772: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5309,
        in1(1) => S5295,
        out1 => S5357
    );
nor_n_5773: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5357,
        in1(1) => S5342,
        out1 => S5358
    );
nand_n_5774: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5358,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S5359
    );
nor_n_5775: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5342,
        in1(1) => S5321,
        out1 => S5360
    );
nand_n_5776: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5341,
        in1(1) => S5320,
        out1 => S5361
    );
nand_n_5777: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5360,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S5362
    );
nor_n_5778: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5335,
        in1(1) => S5321,
        out1 => S5363
    );
nand_n_5779: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5334,
        in1(1) => S5320,
        out1 => S5364
    );
nand_n_5780: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5363,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S5366
    );
nor_n_5781: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5333,
        in1(1) => S5318,
        out1 => S5367
    );
nand_n_5782: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5331,
        in1(1) => S5317,
        out1 => S5368
    );
nand_n_5783: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5367,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S5369
    );
nor_n_5784: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5357,
        in1(1) => S5335,
        out1 => S5370
    );
nand_n_5785: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5370,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S5371
    );
nor_n_5786: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5357,
        in1(1) => S5318,
        out1 => S5372
    );
nand_n_5787: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5356,
        in1(1) => S5317,
        out1 => S5373
    );
nand_n_5788: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5372,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S5374
    );
nor_n_5789: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5357,
        in1(1) => S5327,
        out1 => S5375
    );
nand_n_5790: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5375,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S5377
    );
nand_n_5791: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5369,
        in1(1) => S5325,
        out1 => S5378
    );
nand_n_5792: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5371,
        in1(1) => S5350,
        out1 => S5379
    );
nor_n_5793: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5379,
        in1(1) => S5378,
        out1 => S5380
    );
nand_n_5794: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5377,
        in1(1) => S5355,
        out1 => S5381
    );
nand_n_5795: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5362,
        in1(1) => S5359,
        out1 => S5382
    );
nor_n_5796: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5382,
        in1(1) => S5381,
        out1 => S5383
    );
nand_n_5797: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5383,
        in1(1) => S5380,
        out1 => S5384
    );
nand_n_5798: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5366,
        in1(1) => S5330,
        out1 => S5385
    );
nor_n_5799: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5385,
        in1(1) => S5348,
        out1 => S5386
    );
nand_n_5800: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5374,
        in1(1) => S5352,
        out1 => S5388
    );
nor_n_5801: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5340,
        in1(1) => S5318,
        out1 => S5389
    );
nand_n_5802: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5339,
        in1(1) => S5317,
        out1 => S5390
    );
nor_n_5803: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5390,
        in1(1) => S5966,
        out1 => S5391
    );
nand_n_5804: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5389,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S5392
    );
nand_n_5805: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5392,
        in1(1) => S5338,
        out1 => S5393
    );
nor_n_5806: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5393,
        in1(1) => S5388,
        out1 => S5394
    );
nand_n_5807: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5394,
        in1(1) => S5386,
        out1 => S5395
    );
nor_n_5808: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5342,
        in1(1) => S5333,
        out1 => S5396
    );
nor_n_5809: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5395,
        in1(1) => S5384,
        out1 => S5397
    );
notg_5810: ENTITY WORK.notg
    PORT MAP (
        in1 => S5397,
        out1 => new_datapath_shiftunit_1961_A
    );
nand_n_5811: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5323,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S5399
    );
nand_n_5812: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5363,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S5400
    );
nand_n_5813: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5360,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S5401
    );
nand_n_5814: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5356,
        in1(1) => S5351,
        out1 => S5402
    );
nand_n_5815: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5353,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S5403
    );
nand_n_5816: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5370,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S5404
    );
nand_n_5817: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5349,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S5405
    );
nand_n_5818: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5336,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S5406
    );
notg_5819: ENTITY WORK.notg
    PORT MAP (
        in1 => S5406,
        out1 => S5407
    );
nand_n_5820: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5375,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S5409
    );
nand_n_5821: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5372,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S5410
    );
nand_n_5822: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5367,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S5411
    );
nand_n_5823: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5344,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S5412
    );
notg_5824: ENTITY WORK.notg
    PORT MAP (
        in1 => S5412,
        out1 => S5413
    );
nand_n_5825: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5346,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S5414
    );
nand_n_5826: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5328,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S5415
    );
nand_n_5827: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5414,
        in1(1) => S5410,
        out1 => S5416
    );
nand_n_5828: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5401,
        in1(1) => S5399,
        out1 => S5417
    );
nor_n_5829: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5417,
        in1(1) => S5416,
        out1 => S5418
    );
nor_n_5830: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5390,
        in1(1) => S5957,
        out1 => S5420
    );
nor_n_5831: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S4652,
        in1(1) => S3401,
        out1 => S5421
    );
nand_n_5832: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S4653,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S5422
    );
nor_n_5833: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5422,
        in1(1) => S5315,
        out1 => S5423
    );
nand_n_5834: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5421,
        in1(1) => S5341,
        out1 => S5424
    );
notg_5835: ENTITY WORK.notg
    PORT MAP (
        in1 => S5424,
        out1 => S5425
    );
nor_n_5836: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5424,
        in1(1) => S5333,
        out1 => S5426
    );
nor_n_5837: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5426,
        in1(1) => S5420,
        out1 => S5427
    );
nand_n_5838: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5409,
        in1(1) => S5400,
        out1 => S5428
    );
nor_n_5839: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5428,
        in1(1) => S5407,
        out1 => S5429
    );
nand_n_5840: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5429,
        in1(1) => S5427,
        out1 => S5431
    );
nand_n_5841: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5415,
        in1(1) => S5402,
        out1 => S5432
    );
nor_n_5842: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5432,
        in1(1) => S5413,
        out1 => S5433
    );
nand_n_5843: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5411,
        in1(1) => S5404,
        out1 => S5434
    );
nand_n_5844: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5405,
        in1(1) => S5403,
        out1 => S5435
    );
nor_n_5845: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5435,
        in1(1) => S5434,
        out1 => S5436
    );
nand_n_5846: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5436,
        in1(1) => S5433,
        out1 => S5437
    );
nor_n_5847: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5437,
        in1(1) => S5431,
        out1 => S5438
    );
nand_n_5848: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5438,
        in1(1) => S5418,
        out1 => new_datapath_shiftunit_1979_A
    );
nor_n_5849: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5324,
        in1(1) => S5957,
        out1 => S5439
    );
nand_n_5850: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5323,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S5441
    );
nand_n_5851: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5372,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S5442
    );
nand_n_5852: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5328,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S5443
    );
nand_n_5853: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5375,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S5444
    );
nand_n_5854: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5349,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S5445
    );
nand_n_5855: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5370,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S5446
    );
nand_n_5856: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5360,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S5447
    );
nand_n_5857: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5353,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S5448
    );
nand_n_5858: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5346,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S5449
    );
nand_n_5859: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5336,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S5450
    );
nand_n_5860: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5423,
        in1(1) => S5309,
        out1 => S5452
    );
nand_n_5861: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5367,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S5453
    );
nor_n_5862: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5364,
        in1(1) => S5916,
        out1 => S5454
    );
nand_n_5863: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5363,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S5455
    );
nand_n_5864: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5344,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S5456
    );
nand_n_5865: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5456,
        in1(1) => S5450,
        out1 => S5457
    );
nor_n_5866: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5457,
        in1(1) => S5439,
        out1 => S5458
    );
nand_n_5867: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5453,
        in1(1) => S5445,
        out1 => S5459
    );
nand_n_5868: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5425,
        in1(1) => S5309,
        out1 => S5460
    );
nand_n_5869: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5460,
        in1(1) => S5447,
        out1 => S5461
    );
nor_n_5870: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5461,
        in1(1) => S5459,
        out1 => S5463
    );
nand_n_5871: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5463,
        in1(1) => S5458,
        out1 => S5464
    );
nand_n_5872: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5448,
        in1(1) => S5443,
        out1 => S5465
    );
nand_n_5873: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5389,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S5466
    );
nand_n_5874: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5466,
        in1(1) => S5444,
        out1 => S5467
    );
nor_n_5875: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5467,
        in1(1) => S5465,
        out1 => S5468
    );
nand_n_5876: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5449,
        in1(1) => S5442,
        out1 => S5469
    );
nand_n_5877: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5455,
        in1(1) => S5446,
        out1 => S5470
    );
nor_n_5878: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5470,
        in1(1) => S5469,
        out1 => S5471
    );
nand_n_5879: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5471,
        in1(1) => S5468,
        out1 => S5472
    );
nor_n_5880: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5472,
        in1(1) => S5464,
        out1 => S5474
    );
notg_5881: ENTITY WORK.notg
    PORT MAP (
        in1 => S5474,
        out1 => new_datapath_shiftunit_1997_A
    );
nor_n_5882: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5364,
        in1(1) => S5907,
        out1 => S5475
    );
nand_n_5883: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5363,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S5476
    );
nand_n_5884: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5367,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S5477
    );
nand_n_5885: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5353,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S5478
    );
nand_n_5886: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5336,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S5479
    );
notg_5887: ENTITY WORK.notg
    PORT MAP (
        in1 => S5479,
        out1 => S5480
    );
nor_n_5888: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5324,
        in1(1) => S5947,
        out1 => S5481
    );
nand_n_5889: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5328,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S5482
    );
notg_5890: ENTITY WORK.notg
    PORT MAP (
        in1 => S5482,
        out1 => S5484
    );
nand_n_5891: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5346,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S5485
    );
nand_n_5892: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5370,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S5486
    );
nand_n_5893: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5321,
        in1(1) => S4652,
        out1 => S5487
    );
nand_n_5894: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5487,
        in1(1) => S5351,
        out1 => S5488
    );
nand_n_5895: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5349,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S5489
    );
nand_n_5896: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5372,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S5490
    );
nand_n_5897: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5375,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S5491
    );
nand_n_5898: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5491,
        in1(1) => S5485,
        out1 => S5492
    );
nor_n_5899: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5492,
        in1(1) => S5484,
        out1 => S5493
    );
nand_n_5900: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5493,
        in1(1) => S5488,
        out1 => S5495
    );
nand_n_5901: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5490,
        in1(1) => S5478,
        out1 => S5496
    );
nand_n_5902: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5389,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S5497
    );
nor_n_5903: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5496,
        in1(1) => S5475,
        out1 => S5498
    );
nor_n_5904: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5481,
        in1(1) => S5480,
        out1 => S5499
    );
nand_n_5905: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5497,
        in1(1) => S5477,
        out1 => S5500
    );
nand_n_5906: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5489,
        in1(1) => S5486,
        out1 => S5501
    );
nor_n_5907: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5501,
        in1(1) => S5500,
        out1 => S5502
    );
nand_n_5908: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5502,
        in1(1) => S5499,
        out1 => S5503
    );
nor_n_5909: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5503,
        in1(1) => S5495,
        out1 => S5504
    );
nand_n_5910: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5504,
        in1(1) => S5498,
        out1 => new_datapath_shiftunit_2015_A
    );
nor_n_5911: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5324,
        in1(1) => S5936,
        out1 => S5506
    );
nand_n_5912: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5323,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S5507
    );
nor_n_5913: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5390,
        in1(1) => S5926,
        out1 => S5508
    );
nand_n_5914: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5389,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S5509
    );
nor_n_5915: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5508,
        in1(1) => S5506,
        out1 => S5510
    );
nand_n_5916: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5375,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S5511
    );
nand_n_5917: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5363,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S5512
    );
nand_n_5918: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5349,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S5513
    );
notg_5919: ENTITY WORK.notg
    PORT MAP (
        in1 => S5513,
        out1 => S5514
    );
nand_n_5920: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5370,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S5516
    );
nor_n_5921: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5373,
        in1(1) => S5916,
        out1 => S5517
    );
nand_n_5922: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5328,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S5518
    );
nand_n_5923: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5353,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S5519
    );
nor_n_5924: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5368,
        in1(1) => S5907,
        out1 => S5520
    );
nand_n_5925: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5367,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S5521
    );
nand_n_5926: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5336,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S5522
    );
nand_n_5927: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5346,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S5523
    );
nor_n_5928: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5520,
        in1(1) => S5517,
        out1 => S5524
    );
nand_n_5929: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5522,
        in1(1) => S5511,
        out1 => S5525
    );
nand_n_5930: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5523,
        in1(1) => S5512,
        out1 => S5527
    );
nand_n_5931: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5519,
        in1(1) => S5424,
        out1 => S5528
    );
nor_n_5932: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5528,
        in1(1) => S5527,
        out1 => S5529
    );
notg_5933: ENTITY WORK.notg
    PORT MAP (
        in1 => S5529,
        out1 => S5530
    );
nor_n_5934: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5530,
        in1(1) => S5525,
        out1 => S5531
    );
nand_n_5935: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5524,
        in1(1) => S5510,
        out1 => S5532
    );
nand_n_5936: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5518,
        in1(1) => S5513,
        out1 => S5533
    );
notg_5937: ENTITY WORK.notg
    PORT MAP (
        in1 => S5533,
        out1 => S5534
    );
nand_n_5938: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5534,
        in1(1) => S5516,
        out1 => S5535
    );
nor_n_5939: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5535,
        in1(1) => S5532,
        out1 => S5536
    );
nand_n_5940: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5536,
        in1(1) => S5531,
        out1 => new_datapath_shiftunit_2033_A
    );
nand_n_5941: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5367,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S5538
    );
nand_n_5942: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5349,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S5539
    );
nand_n_5943: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5421,
        in1(1) => S5353,
        out1 => S5540
    );
nand_n_5944: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5323,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S5541
    );
nand_n_5945: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5363,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S5542
    );
nand_n_5946: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5372,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S5543
    );
nand_n_5947: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5328,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S5544
    );
nand_n_5948: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5544,
        in1(1) => S5543,
        out1 => S5545
    );
nand_n_5949: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5370,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S5546
    );
nand_n_5950: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5375,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S5548
    );
nand_n_5951: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5336,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S5549
    );
nand_n_5952: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5346,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S5550
    );
nand_n_5953: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5546,
        in1(1) => S5542,
        out1 => S5551
    );
notg_5954: ENTITY WORK.notg
    PORT MAP (
        in1 => S5551,
        out1 => S5552
    );
nand_n_5955: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5552,
        in1(1) => S5549,
        out1 => S5553
    );
nand_n_5956: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5548,
        in1(1) => S5538,
        out1 => S5554
    );
nor_n_5957: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5554,
        in1(1) => S5545,
        out1 => S5555
    );
notg_5958: ENTITY WORK.notg
    PORT MAP (
        in1 => S5555,
        out1 => S5556
    );
nor_n_5959: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5556,
        in1(1) => S5553,
        out1 => S5557
    );
nand_n_5960: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5539,
        in1(1) => S5424,
        out1 => S5559
    );
nand_n_5961: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5389,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S5560
    );
nand_n_5962: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5560,
        in1(1) => S5550,
        out1 => S5561
    );
nand_n_5963: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5541,
        in1(1) => S5540,
        out1 => S5562
    );
nor_n_5964: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5562,
        in1(1) => S5561,
        out1 => S5563
    );
notg_5965: ENTITY WORK.notg
    PORT MAP (
        in1 => S5563,
        out1 => S5564
    );
nor_n_5966: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5564,
        in1(1) => S5559,
        out1 => S5565
    );
nand_n_5967: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5565,
        in1(1) => S5557,
        out1 => new_datapath_shiftunit_2051_A
    );
nand_n_5968: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5336,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S5566
    );
nand_n_5969: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5349,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S5567
    );
nand_n_5970: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5567,
        in1(1) => S5566,
        out1 => S5569
    );
nand_n_5971: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5323,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S5570
    );
nand_n_5972: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5370,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S5571
    );
nand_n_5973: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5363,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S5572
    );
nand_n_5974: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5452,
        in1(1) => S5424,
        out1 => S5573
    );
nand_n_5975: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5372,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S5574
    );
nand_n_5976: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5328,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S5575
    );
nand_n_5977: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5575,
        in1(1) => S5574,
        out1 => S5576
    );
nand_n_5978: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5367,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S5577
    );
nand_n_5979: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5346,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S5578
    );
nor_n_5980: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5390,
        in1(1) => S5907,
        out1 => S5580
    );
nand_n_5981: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5389,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S5581
    );
nand_n_5982: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5581,
        in1(1) => S5571,
        out1 => S5582
    );
nor_n_5983: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5582,
        in1(1) => S5569,
        out1 => S5583
    );
nand_n_5984: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5578,
        in1(1) => S5570,
        out1 => S5584
    );
nand_n_5985: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5577,
        in1(1) => S5572,
        out1 => S5585
    );
nor_n_5986: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5585,
        in1(1) => S5584,
        out1 => S5586
    );
nor_n_5987: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5576,
        in1(1) => S5573,
        out1 => S5587
    );
nand_n_5988: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5587,
        in1(1) => S5586,
        out1 => S5588
    );
notg_5989: ENTITY WORK.notg
    PORT MAP (
        in1 => S5588,
        out1 => S5589
    );
nand_n_5990: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5589,
        in1(1) => S5583,
        out1 => new_datapath_shiftunit_2069_A
    );
nand_n_5991: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5323,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S5591
    );
nand_n_5992: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5421,
        in1(1) => S5346,
        out1 => S5592
    );
nand_n_5993: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5328,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S5593
    );
nand_n_5994: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5370,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S5594
    );
nand_n_5995: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5372,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S5595
    );
nand_n_5996: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5363,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S5596
    );
nand_n_5997: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5349,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S5597
    );
nand_n_5998: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5336,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S5598
    );
nand_n_5999: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5367,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S5599
    );
nand_n_6000: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5389,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S5601
    );
nand_n_6001: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5601,
        in1(1) => S5594,
        out1 => S5602
    );
nand_n_6002: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5597,
        in1(1) => S5593,
        out1 => S5603
    );
nor_n_6003: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5603,
        in1(1) => S5602,
        out1 => S5604
    );
nand_n_6004: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5595,
        in1(1) => S5592,
        out1 => S5605
    );
nand_n_6005: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5599,
        in1(1) => S5591,
        out1 => S5606
    );
nor_n_6006: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5606,
        in1(1) => S5605,
        out1 => S5607
    );
nand_n_6007: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5598,
        in1(1) => S5596,
        out1 => S5608
    );
nor_n_6008: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5608,
        in1(1) => S5573,
        out1 => S5609
    );
nand_n_6009: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5609,
        in1(1) => S5607,
        out1 => S5610
    );
notg_6010: ENTITY WORK.notg
    PORT MAP (
        in1 => S5610,
        out1 => S5612
    );
nand_n_6011: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5612,
        in1(1) => S5604,
        out1 => new_datapath_shiftunit_2087_A
    );
nand_n_6012: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5349,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S5613
    );
nand_n_6013: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5370,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S5614
    );
nand_n_6014: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5336,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S5615
    );
nand_n_6015: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5323,
        in1(1) => new_datapath_addsubunit_in1_8,
        out1 => S5616
    );
nand_n_6016: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5389,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S5617
    );
nand_n_6017: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5617,
        in1(1) => S5616,
        out1 => S5618
    );
notg_6018: ENTITY WORK.notg
    PORT MAP (
        in1 => S5618,
        out1 => S5619
    );
nor_n_6019: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5368,
        in1(1) => S3357,
        out1 => S5620
    );
nand_n_6020: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5367,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S5622
    );
nor_n_6021: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5620,
        in1(1) => S5423,
        out1 => S5623
    );
nand_n_6022: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5363,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S5624
    );
nand_n_6023: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5372,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S5625
    );
nand_n_6024: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5625,
        in1(1) => S5624,
        out1 => S5626
    );
nand_n_6025: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5614,
        in1(1) => S5613,
        out1 => S5627
    );
nor_n_6026: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5627,
        in1(1) => S5626,
        out1 => S5628
    );
notg_6027: ENTITY WORK.notg
    PORT MAP (
        in1 => S5628,
        out1 => S5629
    );
nand_n_6028: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5619,
        in1(1) => S5615,
        out1 => S5630
    );
nor_n_6029: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5630,
        in1(1) => S5629,
        out1 => S5631
    );
nand_n_6030: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5631,
        in1(1) => S5623,
        out1 => new_datapath_shiftunit_2105_A
    );
nand_n_6031: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5363,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S5633
    );
nand_n_6032: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5372,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S5634
    );
nand_n_6033: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5367,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S5635
    );
nand_n_6034: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5349,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S5636
    );
nor_n_6035: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5370,
        in1(1) => S4653,
        out1 => S5637
    );
nand_n_6036: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5309,
        in1(1) => S5303,
        out1 => S5638
    );
notg_6037: ENTITY WORK.notg
    PORT MAP (
        in1 => S5638,
        out1 => S5639
    );
nor_n_6038: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5639,
        in1(1) => S5316,
        out1 => S5640
    );
nand_n_6039: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5638,
        in1(1) => S5315,
        out1 => S5641
    );
nor_n_6040: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5637,
        in1(1) => S3401,
        out1 => S5643
    );
nand_n_6041: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5643,
        in1(1) => S5641,
        out1 => S5644
    );
nand_n_6042: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5323,
        in1(1) => new_datapath_addsubunit_in1_9,
        out1 => S5645
    );
nand_n_6043: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5645,
        in1(1) => S5644,
        out1 => S5646
    );
nand_n_6044: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5389,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S5647
    );
nand_n_6045: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5635,
        in1(1) => S5633,
        out1 => S5648
    );
nand_n_6046: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5636,
        in1(1) => S5634,
        out1 => S5649
    );
nor_n_6047: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5649,
        in1(1) => S5648,
        out1 => S5650
    );
nand_n_6048: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5650,
        in1(1) => S5647,
        out1 => S5651
    );
nor_n_6049: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5651,
        in1(1) => S5646,
        out1 => S5652
    );
notg_6050: ENTITY WORK.notg
    PORT MAP (
        in1 => S5652,
        out1 => new_datapath_shiftunit_2123_A
    );
nand_n_6051: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5349,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S5654
    );
nand_n_6052: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5363,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S5655
    );
nand_n_6053: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5655,
        in1(1) => S5654,
        out1 => S5656
    );
nand_n_6054: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5372,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S5657
    );
nand_n_6055: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5367,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S5658
    );
nand_n_6056: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5323,
        in1(1) => new_datapath_addsubunit_in1_10,
        out1 => S5659
    );
nor_n_6057: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5640,
        in1(1) => S5422,
        out1 => S5660
    );
nor_n_6058: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5660,
        in1(1) => S5656,
        out1 => S5661
    );
nand_n_6059: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5389,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S5662
    );
nand_n_6060: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5662,
        in1(1) => S5657,
        out1 => S5664
    );
nand_n_6061: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5659,
        in1(1) => S5658,
        out1 => S5665
    );
nor_n_6062: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5665,
        in1(1) => S5664,
        out1 => S5666
    );
nand_n_6063: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5666,
        in1(1) => S5661,
        out1 => new_datapath_shiftunit_2141_A
    );
nand_n_6064: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5421,
        in1(1) => S5349,
        out1 => S5667
    );
nand_n_6065: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5367,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S5668
    );
nand_n_6066: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5668,
        in1(1) => S5667,
        out1 => S5669
    );
nand_n_6067: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5372,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S5670
    );
nand_n_6068: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5363,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S5671
    );
nand_n_6069: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5323,
        in1(1) => new_datapath_addsubunit_in1_11,
        out1 => S5672
    );
nand_n_6070: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5672,
        in1(1) => S5670,
        out1 => S5674
    );
nand_n_6071: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5389,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S5675
    );
nand_n_6072: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5675,
        in1(1) => S5671,
        out1 => S5676
    );
nor_n_6073: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5676,
        in1(1) => S5674,
        out1 => S5677
    );
nor_n_6074: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5669,
        in1(1) => S5660,
        out1 => S5678
    );
nand_n_6075: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5678,
        in1(1) => S5677,
        out1 => new_datapath_shiftunit_2159_A
    );
nand_n_6076: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5323,
        in1(1) => new_datapath_addsubunit_in1_12,
        out1 => S5679
    );
nand_n_6077: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5372,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S5680
    );
nor_n_6078: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5331,
        in1(1) => S5318,
        out1 => S5681
    );
nand_n_6079: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5318,
        in1(1) => S4652,
        out1 => S5682
    );
nand_n_6080: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5682,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S5684
    );
nor_n_6081: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5684,
        in1(1) => S5681,
        out1 => S5685
    );
nand_n_6082: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5389,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S5686
    );
nand_n_6083: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5686,
        in1(1) => S5680,
        out1 => S5687
    );
nor_n_6084: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5687,
        in1(1) => S5685,
        out1 => S5688
    );
nand_n_6085: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5688,
        in1(1) => S5679,
        out1 => new_datapath_shiftunit_2177_A
    );
nor_n_6086: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5681,
        in1(1) => S4652,
        out1 => S5689
    );
nor_n_6087: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5689,
        in1(1) => S5372,
        out1 => S5690
    );
nor_n_6088: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5690,
        in1(1) => S3401,
        out1 => S5691
    );
nand_n_6089: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5323,
        in1(1) => new_datapath_addsubunit_in1_13,
        out1 => S5692
    );
nand_n_6090: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5389,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S5694
    );
nand_n_6091: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5694,
        in1(1) => S5692,
        out1 => S5695
    );
nor_n_6092: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5695,
        in1(1) => S5691,
        out1 => S5696
    );
notg_6093: ENTITY WORK.notg
    PORT MAP (
        in1 => S5696,
        out1 => new_datapath_shiftunit_2195_A
    );
nor_n_6094: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5422,
        in1(1) => S5319,
        out1 => S5697
    );
nand_n_6095: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5323,
        in1(1) => new_datapath_addsubunit_in1_14,
        out1 => S5698
    );
nand_n_6096: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5389,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S5699
    );
notg_6097: ENTITY WORK.notg
    PORT MAP (
        in1 => S5699,
        out1 => S5700
    );
nor_n_6098: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5700,
        in1(1) => S5697,
        out1 => S5701
    );
nand_n_6099: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5701,
        in1(1) => S5698,
        out1 => new_datapath_shiftunit_2213_A
    );
nand_n_6100: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5323,
        in1(1) => new_datapath_addsubunit_in1_15,
        out1 => S5703
    );
nand_n_6101: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5703,
        in1(1) => S5422,
        out1 => new_datapath_shiftunit_2231_A
    );
nand_n_6102: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5389,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S5704
    );
nand_n_6103: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5704,
        in1(1) => S5399,
        out1 => new_datapath_shiftunit_2283_A
    );
nor_n_6104: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5373,
        in1(1) => S5975,
        out1 => S5705
    );
nor_n_6105: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5705,
        in1(1) => S5391,
        out1 => S5706
    );
nand_n_6106: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5706,
        in1(1) => S5441,
        out1 => new_datapath_shiftunit_2301_A
    );
nor_n_6107: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5373,
        in1(1) => S5966,
        out1 => S5707
    );
nor_n_6108: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5368,
        in1(1) => S5975,
        out1 => S5708
    );
nor_n_6109: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5707,
        in1(1) => S5420,
        out1 => S5709
    );
nor_n_6110: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5708,
        in1(1) => S5481,
        out1 => S5711
    );
nand_n_6111: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5711,
        in1(1) => S5709,
        out1 => new_datapath_shiftunit_2319_A
    );
nand_n_6112: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5367,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S5712
    );
nand_n_6113: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5363,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S5713
    );
nand_n_6114: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5712,
        in1(1) => S5507,
        out1 => S5714
    );
nand_n_6115: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5466,
        in1(1) => S5374,
        out1 => S5715
    );
nor_n_6116: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5715,
        in1(1) => S5714,
        out1 => S5716
    );
nand_n_6117: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5716,
        in1(1) => S5713,
        out1 => new_datapath_shiftunit_2337_A
    );
nand_n_6118: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5367,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S5717
    );
nand_n_6119: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5349,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S5718
    );
nand_n_6120: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5718,
        in1(1) => S5717,
        out1 => S5720
    );
notg_6121: ENTITY WORK.notg
    PORT MAP (
        in1 => S5720,
        out1 => S5721
    );
nand_n_6122: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5363,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S5722
    );
nand_n_6123: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5497,
        in1(1) => S5410,
        out1 => S5723
    );
nand_n_6124: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5722,
        in1(1) => S5541,
        out1 => S5724
    );
nor_n_6125: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5724,
        in1(1) => S5723,
        out1 => S5725
    );
nand_n_6126: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5725,
        in1(1) => S5721,
        out1 => new_datapath_shiftunit_2355_A
    );
nor_n_6127: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5364,
        in1(1) => S5957,
        out1 => S5726
    );
nand_n_6128: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5349,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S5727
    );
nand_n_6129: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5370,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S5728
    );
nand_n_6130: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5442,
        in1(1) => S5369,
        out1 => S5730
    );
nand_n_6131: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5727,
        in1(1) => S5509,
        out1 => S5731
    );
nor_n_6132: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5731,
        in1(1) => S5726,
        out1 => S5732
    );
nand_n_6133: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5728,
        in1(1) => S5570,
        out1 => S5733
    );
nor_n_6134: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5733,
        in1(1) => S5730,
        out1 => S5734
    );
nand_n_6135: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5734,
        in1(1) => S5732,
        out1 => new_datapath_shiftunit_2373_A
    );
nand_n_6136: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5490,
        in1(1) => S5411,
        out1 => S5735
    );
nand_n_6137: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5591,
        in1(1) => S5560,
        out1 => S5736
    );
nor_n_6138: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5736,
        in1(1) => S5735,
        out1 => S5737
    );
nand_n_6139: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5370,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S5738
    );
nand_n_6140: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5363,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S5740
    );
nand_n_6141: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5740,
        in1(1) => S5738,
        out1 => S5741
    );
nand_n_6142: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5336,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S5742
    );
nand_n_6143: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5349,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S5743
    );
nand_n_6144: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5743,
        in1(1) => S5742,
        out1 => S5744
    );
nor_n_6145: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5744,
        in1(1) => S5741,
        out1 => S5745
    );
nand_n_6146: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5745,
        in1(1) => S5737,
        out1 => new_datapath_shiftunit_2391_A
    );
nand_n_6147: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5349,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S5746
    );
nand_n_6148: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5370,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S5747
    );
nor_n_6149: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5329,
        in1(1) => S5975,
        out1 => S5748
    );
nand_n_6150: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5336,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S5750
    );
nand_n_6151: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5747,
        in1(1) => S5746,
        out1 => S5751
    );
nor_n_6152: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5580,
        in1(1) => S5517,
        out1 => S5752
    );
nand_n_6153: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5752,
        in1(1) => S5750,
        out1 => S5753
    );
nor_n_6154: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5753,
        in1(1) => S5751,
        out1 => S5754
    );
nand_n_6155: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5616,
        in1(1) => S5453,
        out1 => S5755
    );
notg_6156: ENTITY WORK.notg
    PORT MAP (
        in1 => S5755,
        out1 => S5756
    );
nand_n_6157: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5756,
        in1(1) => S5366,
        out1 => S5757
    );
nor_n_6158: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5757,
        in1(1) => S5748,
        out1 => S5758
    );
nand_n_6159: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5758,
        in1(1) => S5754,
        out1 => new_datapath_shiftunit_2409_A
    );
nand_n_6160: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5370,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S5760
    );
nand_n_6161: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5349,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S5761
    );
nand_n_6162: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5761,
        in1(1) => S5760,
        out1 => S5762
    );
nand_n_6163: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5336,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S5763
    );
nand_n_6164: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5346,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S5764
    );
nand_n_6165: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5764,
        in1(1) => S5763,
        out1 => S5765
    );
nor_n_6166: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5765,
        in1(1) => S5762,
        out1 => S5766
    );
nand_n_6167: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5645,
        in1(1) => S5601,
        out1 => S5767
    );
nand_n_6168: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5477,
        in1(1) => S5400,
        out1 => S5768
    );
nand_n_6169: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5328,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S5769
    );
nand_n_6170: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5769,
        in1(1) => S5543,
        out1 => S5771
    );
nor_n_6171: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5771,
        in1(1) => S5768,
        out1 => S5772
    );
notg_6172: ENTITY WORK.notg
    PORT MAP (
        in1 => S5772,
        out1 => S5773
    );
nor_n_6173: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5773,
        in1(1) => S5767,
        out1 => S5774
    );
nand_n_6174: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5774,
        in1(1) => S5766,
        out1 => new_datapath_shiftunit_2427_A
    );
nand_n_6175: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5336,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S5775
    );
nand_n_6176: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5328,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S5776
    );
nand_n_6177: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5375,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S5777
    );
nand_n_6178: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5346,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S5778
    );
nand_n_6179: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5370,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S5779
    );
nand_n_6180: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5659,
        in1(1) => S5521,
        out1 => S5781
    );
nor_n_6181: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5781,
        in1(1) => S5454,
        out1 => S5782
    );
nand_n_6182: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5617,
        in1(1) => S5574,
        out1 => S5783
    );
nand_n_6183: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5775,
        in1(1) => S5350,
        out1 => S5784
    );
nor_n_6184: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5784,
        in1(1) => S5783,
        out1 => S5785
    );
nand_n_6185: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5785,
        in1(1) => S5782,
        out1 => S5786
    );
notg_6186: ENTITY WORK.notg
    PORT MAP (
        in1 => S5786,
        out1 => S5787
    );
nand_n_6187: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5778,
        in1(1) => S5777,
        out1 => S5788
    );
nand_n_6188: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5779,
        in1(1) => S5776,
        out1 => S5789
    );
nor_n_6189: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5789,
        in1(1) => S5788,
        out1 => S5790
    );
nand_n_6190: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5790,
        in1(1) => S5787,
        out1 => new_datapath_shiftunit_2445_A
    );
nand_n_6191: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5346,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S5792
    );
nand_n_6192: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5328,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S5793
    );
nand_n_6193: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5353,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S5794
    );
nand_n_6194: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5370,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S5795
    );
nand_n_6195: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5375,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S5796
    );
nand_n_6196: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5336,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S5797
    );
nand_n_6197: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5794,
        in1(1) => S5647,
        out1 => S5798
    );
nand_n_6198: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5796,
        in1(1) => S5405,
        out1 => S5799
    );
nor_n_6199: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5799,
        in1(1) => S5798,
        out1 => S5800
    );
notg_6200: ENTITY WORK.notg
    PORT MAP (
        in1 => S5800,
        out1 => S5801
    );
nand_n_6201: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5797,
        in1(1) => S5538,
        out1 => S5802
    );
nor_n_6202: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5802,
        in1(1) => S5801,
        out1 => S5803
    );
nand_n_6203: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5792,
        in1(1) => S5595,
        out1 => S5804
    );
nand_n_6204: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5672,
        in1(1) => S5476,
        out1 => S5805
    );
nand_n_6205: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5795,
        in1(1) => S5793,
        out1 => S5806
    );
nor_n_6206: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5806,
        in1(1) => S5805,
        out1 => S5807
    );
notg_6207: ENTITY WORK.notg
    PORT MAP (
        in1 => S5807,
        out1 => S5808
    );
nor_n_6208: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5808,
        in1(1) => S5804,
        out1 => S5809
    );
nand_n_6209: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5809,
        in1(1) => S5803,
        out1 => new_datapath_shiftunit_2463_A
    );
nand_n_6210: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5679,
        in1(1) => S5662,
        out1 => S5811
    );
nand_n_6211: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5353,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S5812
    );
nand_n_6212: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5328,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S5813
    );
nand_n_6213: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5346,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S5814
    );
nor_n_6214: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5337,
        in1(1) => S5926,
        out1 => S5815
    );
nand_n_6215: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5360,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S5816
    );
nand_n_6216: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5375,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S5817
    );
nand_n_6217: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5512,
        in1(1) => S5445,
        out1 => S5818
    );
nor_n_6218: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5818,
        in1(1) => S5815,
        out1 => S5819
    );
nand_n_6219: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5817,
        in1(1) => S5814,
        out1 => S5820
    );
nand_n_6220: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5816,
        in1(1) => S5813,
        out1 => S5822
    );
nor_n_6221: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5822,
        in1(1) => S5820,
        out1 => S5823
    );
nand_n_6222: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5823,
        in1(1) => S5819,
        out1 => S5824
    );
notg_6223: ENTITY WORK.notg
    PORT MAP (
        in1 => S5824,
        out1 => S5825
    );
nand_n_6224: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5812,
        in1(1) => S5625,
        out1 => S5826
    );
nor_n_6225: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5826,
        in1(1) => S5811,
        out1 => S5827
    );
notg_6226: ENTITY WORK.notg
    PORT MAP (
        in1 => S5827,
        out1 => S5828
    );
nand_n_6227: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5577,
        in1(1) => S5371,
        out1 => S5829
    );
nor_n_6228: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5829,
        in1(1) => S5828,
        out1 => S5830
    );
nand_n_6229: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5830,
        in1(1) => S5825,
        out1 => new_datapath_shiftunit_2481_A
    );
nand_n_6230: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5353,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S5831
    );
nand_n_6231: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5346,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S5832
    );
nand_n_6232: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5360,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S5833
    );
nand_n_6233: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5328,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S5834
    );
nand_n_6234: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5336,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S5835
    );
nand_n_6235: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5344,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S5836
    );
nand_n_6236: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5375,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S5837
    );
nand_n_6237: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5836,
        in1(1) => S5833,
        out1 => S5838
    );
nand_n_6238: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5834,
        in1(1) => S5599,
        out1 => S5839
    );
nor_n_6239: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5839,
        in1(1) => S5838,
        out1 => S5840
    );
notg_6240: ENTITY WORK.notg
    PORT MAP (
        in1 => S5840,
        out1 => S5842
    );
nand_n_6241: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5835,
        in1(1) => S5675,
        out1 => S5843
    );
nor_n_6242: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5843,
        in1(1) => S5842,
        out1 => S5844
    );
nand_n_6243: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5831,
        in1(1) => S5692,
        out1 => S5845
    );
nand_n_6244: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5542,
        in1(1) => S5489,
        out1 => S5846
    );
nor_n_6245: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5846,
        in1(1) => S5845,
        out1 => S5847
    );
nand_n_6246: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5837,
        in1(1) => S5404,
        out1 => S5848
    );
nand_n_6247: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5832,
        in1(1) => S5634,
        out1 => S5849
    );
nor_n_6248: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5849,
        in1(1) => S5848,
        out1 => S5850
    );
nand_n_6249: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5850,
        in1(1) => S5847,
        out1 => S5851
    );
notg_6250: ENTITY WORK.notg
    PORT MAP (
        in1 => S5851,
        out1 => S5853
    );
nand_n_6251: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5853,
        in1(1) => S5844,
        out1 => new_datapath_shiftunit_2499_A
    );
nand_n_6252: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5446,
        in1(1) => S5338,
        out1 => S5854
    );
nand_n_6253: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5360,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S5855
    );
nand_n_6254: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5358,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S5856
    );
nand_n_6255: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5375,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S5857
    );
nand_n_6256: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5344,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S5858
    );
nand_n_6257: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5353,
        in1(1) => new_datapath_addsubunit_in1_3,
        out1 => S5859
    );
nand_n_6258: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5328,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S5860
    );
nand_n_6259: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5346,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S5861
    );
nand_n_6260: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5657,
        in1(1) => S5622,
        out1 => S5863
    );
nor_n_6261: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5863,
        in1(1) => S5854,
        out1 => S5864
    );
nand_n_6262: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5861,
        in1(1) => S5857,
        out1 => S5865
    );
nand_n_6263: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5859,
        in1(1) => S5855,
        out1 => S5866
    );
nor_n_6264: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5866,
        in1(1) => S5865,
        out1 => S5867
    );
nand_n_6265: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5867,
        in1(1) => S5864,
        out1 => S5868
    );
nand_n_6266: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5860,
        in1(1) => S5856,
        out1 => S5869
    );
nand_n_6267: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5858,
        in1(1) => S5698,
        out1 => S5870
    );
nor_n_6268: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5870,
        in1(1) => S5869,
        out1 => S5871
    );
nand_n_6269: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5686,
        in1(1) => S5572,
        out1 => S5872
    );
nor_n_6270: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5872,
        in1(1) => S5514,
        out1 => S5873
    );
nand_n_6271: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5873,
        in1(1) => S5871,
        out1 => S5874
    );
nor_n_6272: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5874,
        in1(1) => S5868,
        out1 => S5875
    );
notg_6273: ENTITY WORK.notg
    PORT MAP (
        in1 => S5875,
        out1 => new_datapath_shiftunit_2517_A
    );
nor_n_6274: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5361,
        in1(1) => S5947,
        out1 => S5876
    );
nand_n_6275: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5358,
        in1(1) => new_datapath_addsubunit_in1_1,
        out1 => S5877
    );
nand_n_6276: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5396,
        in1(1) => new_datapath_addsubunit_in1_0,
        out1 => S5878
    );
nand_n_6277: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5328,
        in1(1) => new_datapath_addsubunit_in1_7,
        out1 => S5879
    );
nand_n_6278: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5375,
        in1(1) => new_datapath_addsubunit_in1_5,
        out1 => S5880
    );
notg_6279: ENTITY WORK.notg
    PORT MAP (
        in1 => S5880,
        out1 => S5881
    );
nand_n_6280: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5346,
        in1(1) => new_datapath_addsubunit_in1_6,
        out1 => S5883
    );
nand_n_6281: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5344,
        in1(1) => new_datapath_addsubunit_in1_2,
        out1 => S5884
    );
nand_n_6282: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5353,
        in1(1) => new_datapath_addsubunit_in1_4,
        out1 => S5885
    );
nand_n_6283: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5884,
        in1(1) => S5596,
        out1 => S5886
    );
nor_n_6284: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5886,
        in1(1) => S5876,
        out1 => S5887
    );
nand_n_6285: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5887,
        in1(1) => S5878,
        out1 => S5888
    );
nand_n_6286: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5635,
        in1(1) => S5406,
        out1 => S5889
    );
nor_n_6287: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5889,
        in1(1) => S5888,
        out1 => S5890
    );
nand_n_6288: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5670,
        in1(1) => S5539,
        out1 => S5891
    );
notg_6289: ENTITY WORK.notg
    PORT MAP (
        in1 => S5891,
        out1 => S5892
    );
nand_n_6290: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5892,
        in1(1) => S5877,
        out1 => S5894
    );
nand_n_6291: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5883,
        in1(1) => S5879,
        out1 => S5895
    );
nor_n_6292: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5895,
        in1(1) => S5881,
        out1 => S5896
    );
nand_n_6293: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5703,
        in1(1) => S5486,
        out1 => S5897
    );
nand_n_6294: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5885,
        in1(1) => S5694,
        out1 => S5898
    );
nor_n_6295: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5898,
        in1(1) => S5897,
        out1 => S5899
    );
nand_n_6296: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5899,
        in1(1) => S5896,
        out1 => S5900
    );
nor_n_6297: ENTITY WORK.nor_n
    PORT MAP (
        in1(0) => S5900,
        in1(1) => S5894,
        out1 => S5901
    );
nand_n_6298: ENTITY WORK.nand_n
    PORT MAP (
        in1(0) => S5901,
        in1(1) => S5890,
        out1 => new_datapath_shiftunit_2534_A
    );
bufg_6299: ENTITY WORK.bufg
    PORT MAP (
        in1 => new_controller_outflag_7,
        out1 => S3
    );
bufg_6300: ENTITY WORK.bufg
    PORT MAP (
        in1 => new_controller_outflag_0,
        out1 => S66
    );
bufg_6301: ENTITY WORK.bufg
    PORT MAP (
        in1 => new_controller_outflag_1,
        out1 => S67
    );
bufg_6302: ENTITY WORK.bufg
    PORT MAP (
        in1 => new_controller_outflag_2,
        out1 => S68
    );
bufg_6303: ENTITY WORK.bufg
    PORT MAP (
        in1 => new_controller_outflag_3,
        out1 => S69
    );
bufg_6304: ENTITY WORK.bufg
    PORT MAP (
        in1 => new_controller_outflag_6,
        out1 => S72
    );
dff_6305: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => new_controller_1423_Y_0,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_pstate_0,
        Si => Si_3_sig,
        global_reset => '0'
    );
dff_6306: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => new_controller_1423_Y_1,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_pstate_1,
        Si => new_controller_pstate_0,
        global_reset => '0'
    );
dff_6307: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S73,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_adr_outreg_0,
        Si => new_controller_pstate_1,
        global_reset => '0'
    );
dff_6308: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S74,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_adr_outreg_1,
        Si => new_datapath_adr_outreg_0,
        global_reset => '0'
    );
dff_6309: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S75,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_adr_outreg_2,
        Si => new_datapath_adr_outreg_1,
        global_reset => '0'
    );
dff_6310: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S76,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_adr_outreg_3,
        Si => new_datapath_adr_outreg_2,
        global_reset => '0'
    );
dff_6311: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S77,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_adr_outreg_4,
        Si => new_datapath_adr_outreg_3,
        global_reset => '0'
    );
dff_6312: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S78,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_adr_outreg_5,
        Si => new_datapath_adr_outreg_4,
        global_reset => '0'
    );
dff_6313: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S79,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_adr_outreg_6,
        Si => new_datapath_adr_outreg_5,
        global_reset => '0'
    );

dff_6314: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S80,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_adr_outreg_7,
        Si => new_datapath_adr_outreg_6,
        global_reset => '0'
    );
dff_6315: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S81,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_adr_outreg_8,
        Si => new_datapath_adr_outreg_7,
        global_reset => '0'
    );
dff_6316: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S82,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_adr_outreg_9,
        Si => new_datapath_adr_outreg_8,
        global_reset => '0'
    );
dff_6317: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S83,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_adr_outreg_10,
        Si => new_datapath_adr_outreg_9,
        global_reset => '0'
    );
dff_6318: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S84,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_adr_outreg_11,
        Si => new_datapath_adr_outreg_10,
        global_reset => '0'
    );
dff_6319: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S85,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_adr_outreg_12,
        Si => new_datapath_adr_outreg_11,
        global_reset => '0'
    );
dff_6320: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S86,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_adr_outreg_13,
        Si => new_datapath_adr_outreg_12,
        global_reset => '0'
    );
dff_6321: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S87,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_adr_outreg_14,
        Si => new_datapath_adr_outreg_13,
        global_reset => '0'
    );
dff_6322: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S4,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_adr_outreg_15,
        Si => new_datapath_adr_outreg_14,
        global_reset => '0'
    );
dff_6323: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S66,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_outflag_0,
        Si => new_datapath_adr_outreg_15,
        global_reset => '0'
    );
dff_6324: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S67,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_outflag_1,
        Si => new_controller_outflag_0,
        global_reset => '0'
    );
dff_6325: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S68,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_outflag_2,
        Si => new_controller_outflag_1,
        global_reset => '0'
    );
dff_6326: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S69,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_outflag_3,
        Si => new_controller_outflag_2,
        global_reset => '0'
    );
dff_6327: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S70,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_407_B_0,
        Si => new_controller_outflag_3,
        global_reset => '0'
    );
dff_6328: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S71,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_407_B_2,
        Si => new_controller_407_B_0,
        global_reset => '0'
    );
dff_6329: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S72,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_outflag_6,
        Si => new_controller_407_B_2,
        global_reset => '0'
    );

So_1_sig <= new_controller_outflag_6; 	-- added for scan insertion

dff_6330: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S3,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_outflag_7,
        Si => Si_4_sig,
        global_reset => '0'
    );
dff_6331: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S51,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_instruction_0,
        Si => new_controller_outflag_7,
        global_reset => '0'
    );
dff_6332: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S52,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_instruction_1,
        Si => new_datapath_instruction_0,
        global_reset => '0'
    );
dff_6333: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S53,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_instruction_2,
        Si => new_datapath_instruction_1,
        global_reset => '0'
    );
dff_6334: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S54,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_instruction_3,
        Si => new_datapath_instruction_2,
        global_reset => '0'
    );
dff_6335: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S55,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_fib_0,
        Si => new_datapath_instruction_3,
        global_reset => '0'
    );
dff_6336: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S56,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_fib_1,
        Si => new_controller_fib_0,
        global_reset => '0'
    );
dff_6337: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S57,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_fib_2,
        Si => new_controller_fib_1,
        global_reset => '0'
    );
dff_6338: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S58,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_fib_3,
        Si => new_controller_fib_2,
        global_reset => '0'
    );
dff_6339: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S59,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_fib_4,
        Si => new_controller_fib_3,
        global_reset => '0'
    );
dff_6340: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S60,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_234_B_0,
        Si => new_controller_fib_4,
        global_reset => '0'
    );
dff_6341: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S61,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_opcode_2,
        Si => new_controller_234_B_0,
        global_reset => '0'
    );
dff_6342: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S62,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_opcode_3,
        Si => new_controller_opcode_2,
        global_reset => '0'
    );

dff_6343: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S63,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_opcode_4,
        Si => new_controller_opcode_3,
        global_reset => '0'
    );
dff_6344: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S64,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_opcode_5,
        Si => new_controller_opcode_4,
        global_reset => '0'
    );
dff_6345: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S65,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_opcode_6,
        Si => new_controller_opcode_5,
        global_reset => '0'
    );
dff_6346: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S2,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_controller_opcode_7,
        Si => new_controller_opcode_6,
        global_reset => '0'
    );
dff_6347: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S20,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu1_0,
        Si => new_controller_opcode_7,
        global_reset => '0'
    );
dff_6348: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S21,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu1_1,
        Si => new_datapath_multdivunit_outmdu1_0,
        global_reset => '0'
    );
dff_6349: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S22,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu1_2,
        Si => new_datapath_multdivunit_outmdu1_1,
        global_reset => '0'
    );
dff_6350: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S23,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu1_3,
        Si => new_datapath_multdivunit_outmdu1_2,
        global_reset => '0'
    );
dff_6351: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S24,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu1_4,
        Si => new_datapath_multdivunit_outmdu1_3,
        global_reset => '0'
    );
dff_6352: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S25,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu1_5,
        Si => new_datapath_multdivunit_outmdu1_4,
        global_reset => '0'
    );
dff_6353: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S26,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu1_6,
        Si => new_datapath_multdivunit_outmdu1_5,
        global_reset => '0'
    );
dff_6354: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S27,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu1_7,
        Si => new_datapath_multdivunit_outmdu1_6,
        global_reset => '0'
    );

So_2_sig <= new_datapath_multdivunit_outmdu1_7; 	-- added for scan insertion

dff_6355: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S28,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu1_8,
        Si => Si_5_sig,
        global_reset => '0'
    );
dff_6356: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S29,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu1_9,
        Si => new_datapath_multdivunit_outmdu1_8,
        global_reset => '0'
    );
dff_6357: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S30,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu1_10,
        Si => new_datapath_multdivunit_outmdu1_9,
        global_reset => '0'
    );
dff_6358: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S31,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu1_11,
        Si => new_datapath_multdivunit_outmdu1_10,
        global_reset => '0'
    );
dff_6359: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S32,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu1_12,
        Si => new_datapath_multdivunit_outmdu1_11,
        global_reset => '0'
    );
dff_6360: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S33,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu1_13,
        Si => new_datapath_multdivunit_outmdu1_12,
        global_reset => '0'
    );
dff_6361: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S34,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu1_14,
        Si => new_datapath_multdivunit_outmdu1_13,
        global_reset => '0'
    );
dff_6362: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S35,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu1_15,
        Si => new_datapath_multdivunit_outmdu1_14,
        global_reset => '0'
    );
dff_6363: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S36,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu2_0,
        Si => new_datapath_multdivunit_outmdu1_15,
        global_reset => '0'
    );
dff_6364: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S37,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu2_1,
        Si => new_datapath_multdivunit_outmdu2_0,
        global_reset => '0'
    );
dff_6365: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S38,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu2_2,
        Si => new_datapath_multdivunit_outmdu2_1,
        global_reset => '0'
    );
dff_6366: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S39,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu2_3,
        Si => new_datapath_multdivunit_outmdu2_2,
        global_reset => '0'
    );
dff_6367: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S40,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu2_4,
        Si => new_datapath_multdivunit_outmdu2_3,
        global_reset => '0'
    );
dff_6368: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S41,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu2_5,
        Si => new_datapath_multdivunit_outmdu2_4,
        global_reset => '0'
    );
dff_6369: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S42,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu2_6,
        Si => new_datapath_multdivunit_outmdu2_5,
        global_reset => '0'
    );
dff_6370: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S43,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu2_7,
        Si => new_datapath_multdivunit_outmdu2_6,
        global_reset => '0'
    );
dff_6371: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S44,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu2_8,
        Si => new_datapath_multdivunit_outmdu2_7,
        global_reset => '0'
    );
dff_6372: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S45,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu2_9,
        Si => new_datapath_multdivunit_outmdu2_8,
        global_reset => '0'
    );
dff_6373: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S46,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu2_10,
        Si => new_datapath_multdivunit_outmdu2_9,
        global_reset => '0'
    );
dff_6374: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S47,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu2_11,
        Si => new_datapath_multdivunit_outmdu2_10,
        global_reset => '0'
    );
dff_6375: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S48,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu2_12,
        Si => new_datapath_multdivunit_outmdu2_11,
        global_reset => '0'
    );
dff_6376: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S49,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu2_13,
        Si => new_datapath_multdivunit_outmdu2_12,
        global_reset => '0'
    );
dff_6377: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S50,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu2_14,
        Si => new_datapath_multdivunit_outmdu2_13,
        global_reset => '0'
    );
dff_6378: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S1,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_multdivunit_outmdu2_15,
        Si => new_datapath_multdivunit_outmdu2_14,
        global_reset => '0'
    );
dff_6379: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S5,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_muxmem_in2_0,
        Si => new_datapath_multdivunit_outmdu2_15,
        global_reset => '0'
    );

So_3_sig <= new_datapath_muxmem_in2_0; 	-- added for scan insertion

dff_6380: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S6,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_muxmem_in2_1,
        Si => Si_6_sig,
        global_reset => '0'
    );
dff_6381: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S7,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_muxmem_in2_2,
        Si => new_datapath_muxmem_in2_1,
        global_reset => '0'
    );
dff_6382: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S8,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_muxmem_in2_3,
        Si => new_datapath_muxmem_in2_2,
        global_reset => '0'
    );
dff_6383: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S9,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_muxmem_in2_4,
        Si => new_datapath_muxmem_in2_3,
        global_reset => '0'
    );
dff_6384: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S10,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_muxmem_in2_5,
        Si => new_datapath_muxmem_in2_4,
        global_reset => '0'
    );
dff_6385: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S11,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_muxmem_in2_6,
        Si => new_datapath_muxmem_in2_5,
        global_reset => '0'
    );
dff_6386: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S12,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_muxmem_in2_7,
        Si => new_datapath_muxmem_in2_6,
        global_reset => '0'
    );
dff_6387: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S13,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_muxmem_in2_8,
        Si => new_datapath_muxmem_in2_7,
        global_reset => '0'
    );
dff_6388: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S14,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_muxmem_in2_9,
        Si => new_datapath_muxmem_in2_8,
        global_reset => '0'
    );
dff_6389: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S15,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_muxmem_in2_10,
        Si => new_datapath_muxmem_in2_9,
        global_reset => '0'
    );
dff_6390: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S16,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_muxmem_in2_11,
        Si => new_datapath_muxmem_in2_10,
        global_reset => '0'
    );
dff_6391: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S17,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_muxmem_in2_12,
        Si => new_datapath_muxmem_in2_11,
        global_reset => '0'
    );
dff_6392: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S18,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_muxmem_in2_13,
        Si => new_datapath_muxmem_in2_12,
        global_reset => '0'
    );
dff_6393: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S19,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_muxmem_in2_14,
        Si => new_datapath_muxmem_in2_13,
        global_reset => '0'
    );
dff_6394: ENTITY WORK.dff
    PORT MAP (
        C => new_controller_clk,
        CE => '1',
        CLR => new_controller_rst,
        D => S0,
        NbarT => PbarS_sig,
        PRE => '0',
        Q => new_datapath_muxmem_in2_15,
        Si => new_datapath_muxmem_in2_14,
        global_reset => '0'
    );

fakeDFF_91to100: ENTITY WORK.dffBlock GENERIC MAP (10) 
    PORT MAP (              
        C => new_controller_clk,      	    -- added for scan insertion      
        CE => '0',                 	        -- added for scan insertion         
        CLR => new_controller_rst,      	-- added for scan insertion    
        D => (OTHERS=>'0'),           	    -- added for scan insertion      
        NbarT => PbarS_sig, 	            -- added for scan insertion
        PRE => '0', 	                    -- added for scan insertion
        Q => fakeDFF_sig(9 DOWNTO 0),	    -- added for scan insertion
        Si => new_datapath_muxmem_in2_15,	-- added for scan insertion
        global_reset => '0' 	            -- added for scan insertion
    );

So_4_sig <= fakeDFF_sig(0); 	            -- added for scan insertion
	
pout_6395: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addrbus_0,
        out1 => addrBus(0)
    );
pout_6396: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addrbus_1,
        out1 => addrBus(1)
    );
pout_6397: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addrbus_10,
        out1 => addrBus(10)
    );
pout_6398: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addrbus_11,
        out1 => addrBus(11)
    );
pout_6399: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addrbus_12,
        out1 => addrBus(12)
    );
pout_6400: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addrbus_13,
        out1 => addrBus(13)
    );
pout_6401: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addrbus_14,
        out1 => addrBus(14)
    );
pout_6402: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addrbus_15,
        out1 => addrBus(15)
    );
pout_6403: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addrbus_2,
        out1 => addrBus(2)
    );
pout_6404: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addrbus_3,
        out1 => addrBus(3)
    );
pout_6405: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addrbus_4,
        out1 => addrBus(4)
    );
pout_6406: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addrbus_5,
        out1 => addrBus(5)
    );
pout_6407: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addrbus_6,
        out1 => addrBus(6)
    );
pout_6408: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addrbus_7,
        out1 => addrBus(7)
    );
pout_6409: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addrbus_8,
        out1 => addrBus(8)
    );
pout_6410: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addrbus_9,
        out1 => addrBus(9)
    );
pin_6411: ENTITY WORK.pin
    PORT MAP (
        in1 => clk,
        out1 => new_controller_clk
    );
pin_6412: ENTITY WORK.pin
    PORT MAP (
        in1 => dataBusIn(0),
        out1 => new_datapath_databusin_0
    );
pin_6413: ENTITY WORK.pin
    PORT MAP (
        in1 => dataBusIn(1),
        out1 => new_datapath_databusin_1
    );
pin_6414: ENTITY WORK.pin
    PORT MAP (
        in1 => dataBusIn(10),
        out1 => new_datapath_databusin_10
    );
pin_6415: ENTITY WORK.pin
    PORT MAP (
        in1 => dataBusIn(11),
        out1 => new_datapath_databusin_11
    );
pin_6416: ENTITY WORK.pin
    PORT MAP (
        in1 => dataBusIn(12),
        out1 => new_datapath_databusin_12
    );
pin_6417: ENTITY WORK.pin
    PORT MAP (
        in1 => dataBusIn(13),
        out1 => new_datapath_databusin_13
    );
pin_6418: ENTITY WORK.pin
    PORT MAP (
        in1 => dataBusIn(14),
        out1 => new_datapath_databusin_14
    );
pin_6419: ENTITY WORK.pin
    PORT MAP (
        in1 => dataBusIn(15),
        out1 => new_datapath_databusin_15
    );
pin_6420: ENTITY WORK.pin
    PORT MAP (
        in1 => dataBusIn(2),
        out1 => new_datapath_databusin_2
    );
pin_6421: ENTITY WORK.pin
    PORT MAP (
        in1 => dataBusIn(3),
        out1 => new_datapath_databusin_3
    );
pin_6422: ENTITY WORK.pin
    PORT MAP (
        in1 => dataBusIn(4),
        out1 => new_datapath_databusin_4
    );
pin_6423: ENTITY WORK.pin
    PORT MAP (
        in1 => dataBusIn(5),
        out1 => new_datapath_databusin_5
    );
pin_6424: ENTITY WORK.pin
    PORT MAP (
        in1 => dataBusIn(6),
        out1 => new_datapath_databusin_6
    );
pin_6425: ENTITY WORK.pin
    PORT MAP (
        in1 => dataBusIn(7),
        out1 => new_datapath_databusin_7
    );
pin_6426: ENTITY WORK.pin
    PORT MAP (
        in1 => dataBusIn(8),
        out1 => new_datapath_databusin_8
    );
pin_6427: ENTITY WORK.pin
    PORT MAP (
        in1 => dataBusIn(9),
        out1 => new_datapath_databusin_9
    );
pout_6428: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_0,
        out1 => dataBusOut(0)
    );
pout_6429: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_1,
        out1 => dataBusOut(1)
    );
pout_6430: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_10,
        out1 => dataBusOut(10)
    );
pout_6431: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_11,
        out1 => dataBusOut(11)
    );
pout_6432: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_12,
        out1 => dataBusOut(12)
    );
pout_6433: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_13,
        out1 => dataBusOut(13)
    );
pout_6434: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_14,
        out1 => dataBusOut(14)
    );
pout_6435: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_15,
        out1 => dataBusOut(15)
    );
pout_6436: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_2,
        out1 => dataBusOut(2)
    );
pout_6437: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_3,
        out1 => dataBusOut(3)
    );
pout_6438: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_4,
        out1 => dataBusOut(4)
    );
pout_6439: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_5,
        out1 => dataBusOut(5)
    );
pout_6440: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_6,
        out1 => dataBusOut(6)
    );
pout_6441: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_7,
        out1 => dataBusOut(7)
    );
pout_6442: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_8,
        out1 => dataBusOut(8)
    );
pout_6443: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_addsubunit_in1_9,
        out1 => dataBusOut(9)
    );
pout_6444: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_indatatrf_0,
        out1 => inDataTRF(0)
    );
pout_6445: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_indatatrf_1,
        out1 => inDataTRF(1)
    );
pout_6446: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_indatatrf_10,
        out1 => inDataTRF(10)
    );
pout_6447: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_indatatrf_11,
        out1 => inDataTRF(11)
    );
pout_6448: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_indatatrf_12,
        out1 => inDataTRF(12)
    );
pout_6449: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_indatatrf_13,
        out1 => inDataTRF(13)
    );
pout_6450: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_indatatrf_14,
        out1 => inDataTRF(14)
    );
pout_6451: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_indatatrf_15,
        out1 => inDataTRF(15)
    );
pout_6452: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_indatatrf_2,
        out1 => inDataTRF(2)
    );
pout_6453: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_indatatrf_3,
        out1 => inDataTRF(3)
    );
pout_6454: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_indatatrf_4,
        out1 => inDataTRF(4)
    );
pout_6455: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_indatatrf_5,
        out1 => inDataTRF(5)
    );
pout_6456: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_indatatrf_6,
        out1 => inDataTRF(6)
    );
pout_6457: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_indatatrf_7,
        out1 => inDataTRF(7)
    );
pout_6458: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_indatatrf_8,
        out1 => inDataTRF(8)
    );
pout_6459: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_indatatrf_9,
        out1 => inDataTRF(9)
    );
pout_6460: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_muxrd_outmux_0,
        out1 => outMuxrd(0)
    );
pout_6461: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_muxrd_outmux_1,
        out1 => outMuxrd(1)
    );
pout_6462: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_muxrd_outmux_2,
        out1 => outMuxrd(2)
    );
pout_6463: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_muxrd_outmux_3,
        out1 => outMuxrd(3)
    );
pout_6464: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_muxrs1_outmux_0,
        out1 => outMuxrs1(0)
    );
pout_6465: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_muxrs1_outmux_1,
        out1 => outMuxrs1(1)
    );
pout_6466: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_muxrs1_outmux_2,
        out1 => outMuxrs1(2)
    );
pout_6467: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_muxrs1_outmux_3,
        out1 => outMuxrs1(3)
    );
pout_6468: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_muxrs2_outmux_0,
        out1 => outMuxrs2(0)
    );
pout_6469: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_muxrs2_outmux_1,
        out1 => outMuxrs2(1)
    );
pout_6470: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_muxrs2_outmux_2,
        out1 => outMuxrs2(2)
    );
pout_6471: ENTITY WORK.pout
    PORT MAP (
        in1 => new_datapath_muxrs2_outmux_3,
        out1 => outMuxrs2(3)
    );
pin_6472: ENTITY WORK.pin
    PORT MAP (
        in1 => p1TRF(0),
        out1 => new_datapath_p1trf_0
    );
pin_6473: ENTITY WORK.pin
    PORT MAP (
        in1 => p1TRF(1),
        out1 => new_datapath_p1trf_1
    );
pin_6474: ENTITY WORK.pin
    PORT MAP (
        in1 => p1TRF(10),
        out1 => new_datapath_addsubunit_in1_10
    );
pin_6475: ENTITY WORK.pin
    PORT MAP (
        in1 => p1TRF(11),
        out1 => new_datapath_addsubunit_in1_11
    );
pin_6476: ENTITY WORK.pin
    PORT MAP (
        in1 => p1TRF(12),
        out1 => new_datapath_addsubunit_in1_12
    );
pin_6477: ENTITY WORK.pin
    PORT MAP (
        in1 => p1TRF(13),
        out1 => new_datapath_addsubunit_in1_13
    );
pin_6478: ENTITY WORK.pin
    PORT MAP (
        in1 => p1TRF(14),
        out1 => new_datapath_addsubunit_in1_14
    );
pin_6479: ENTITY WORK.pin
    PORT MAP (
        in1 => p1TRF(15),
        out1 => new_datapath_addsubunit_in1_15
    );
pin_6480: ENTITY WORK.pin
    PORT MAP (
        in1 => p1TRF(2),
        out1 => new_datapath_p1trf_2
    );
pin_6481: ENTITY WORK.pin
    PORT MAP (
        in1 => p1TRF(3),
        out1 => new_datapath_p1trf_3
    );
pin_6482: ENTITY WORK.pin
    PORT MAP (
        in1 => p1TRF(4),
        out1 => new_datapath_p1trf_4
    );
pin_6483: ENTITY WORK.pin
    PORT MAP (
        in1 => p1TRF(5),
        out1 => new_datapath_p1trf_5
    );
pin_6484: ENTITY WORK.pin
    PORT MAP (
        in1 => p1TRF(6),
        out1 => new_datapath_p1trf_6
    );
pin_6485: ENTITY WORK.pin
    PORT MAP (
        in1 => p1TRF(7),
        out1 => new_datapath_p1trf_7
    );
pin_6486: ENTITY WORK.pin
    PORT MAP (
        in1 => p1TRF(8),
        out1 => new_datapath_addsubunit_in1_8
    );
pin_6487: ENTITY WORK.pin
    PORT MAP (
        in1 => p1TRF(9),
        out1 => new_datapath_addsubunit_in1_9
    );
pin_6488: ENTITY WORK.pin
    PORT MAP (
        in1 => p2TRF(0),
        out1 => new_datapath_p2trf_0
    );
pin_6489: ENTITY WORK.pin
    PORT MAP (
        in1 => p2TRF(1),
        out1 => new_datapath_p2trf_1
    );
pin_6490: ENTITY WORK.pin
    PORT MAP (
        in1 => p2TRF(10),
        out1 => new_datapath_multdivunit_1697_B_10
    );
pin_6491: ENTITY WORK.pin
    PORT MAP (
        in1 => p2TRF(11),
        out1 => new_datapath_multdivunit_1697_B_11
    );
pin_6492: ENTITY WORK.pin
    PORT MAP (
        in1 => p2TRF(12),
        out1 => new_datapath_multdivunit_1697_B_12
    );
pin_6493: ENTITY WORK.pin
    PORT MAP (
        in1 => p2TRF(13),
        out1 => new_datapath_multdivunit_1697_B_13
    );
pin_6494: ENTITY WORK.pin
    PORT MAP (
        in1 => p2TRF(14),
        out1 => new_datapath_multdivunit_1697_B_14
    );
pin_6495: ENTITY WORK.pin
    PORT MAP (
        in1 => p2TRF(15),
        out1 => new_datapath_multdivunit_1697_B_15
    );
pin_6496: ENTITY WORK.pin
    PORT MAP (
        in1 => p2TRF(2),
        out1 => new_datapath_p2trf_2
    );
pin_6497: ENTITY WORK.pin
    PORT MAP (
        in1 => p2TRF(3),
        out1 => new_datapath_p2trf_3
    );
pin_6498: ENTITY WORK.pin
    PORT MAP (
        in1 => p2TRF(4),
        out1 => new_datapath_p2trf_4
    );
pin_6499: ENTITY WORK.pin
    PORT MAP (
        in1 => p2TRF(5),
        out1 => new_datapath_p2trf_5
    );
pin_6500: ENTITY WORK.pin
    PORT MAP (
        in1 => p2TRF(6),
        out1 => new_datapath_p2trf_6
    );
pin_6501: ENTITY WORK.pin
    PORT MAP (
        in1 => p2TRF(7),
        out1 => new_datapath_p2trf_7
    );
pin_6502: ENTITY WORK.pin
    PORT MAP (
        in1 => p2TRF(8),
        out1 => new_datapath_multdivunit_1697_B_8
    );
pin_6503: ENTITY WORK.pin
    PORT MAP (
        in1 => p2TRF(9),
        out1 => new_datapath_multdivunit_1697_B_9
    );
pout_6504: ENTITY WORK.pout
    PORT MAP (
        in1 => new_controller_1133_S_0,
        out1 => readInst
    );
pout_6505: ENTITY WORK.pout
    PORT MAP (
        in1 => S6215,
        out1 => readMM
    );
pin_6506: ENTITY WORK.pin
    PORT MAP (
        in1 => readyMEM,
        out1 => new_controller_readymem
    );
pin_6507: ENTITY WORK.pin
    PORT MAP (
        in1 => rst,
        out1 => new_controller_rst
    );
pout_6508: ENTITY WORK.pout
    PORT MAP (
        in1 => S6216,
        out1 => writeMM
    );
pout_6509: ENTITY WORK.pout
    PORT MAP (
        in1 => new_controller_1133_Y,
        out1 => writeTRF
    );
pin_6510: ENTITY WORK.pin               -- added for test insertion
    PORT MAP (                          -- added for test insertion
        in1 => PbarS,                   -- added for test insertion
        out1 => PbarS_sig               -- added for test insertion
    );                                  -- added for test insertion
pin_6511: ENTITY WORK.pin               -- added for test insertion
    PORT MAP (                          -- added for test insertion
        in1 => Si_3,                    -- added for test insertion
        out1 => Si_3_sig                -- added for test insertion
    );                                  -- added for test insertion
pin_6512: ENTITY WORK.pin               -- added for test insertion
    PORT MAP (                          -- added for test insertion
        in1 => Si_4,                    -- added for test insertion
        out1 => Si_4_sig                -- added for test insertion
    );                                  -- added for test insertion
pin_6513: ENTITY WORK.pin               -- added for test insertion
    PORT MAP (                          -- added for test insertion
        in1 => Si_5,                    -- added for test insertion
        out1 => Si_5_sig                -- added for test insertion
    );                                  -- added for test insertion
pin_6514: ENTITY WORK.pin               -- added for test insertion
    PORT MAP (                          -- added for test insertion
        in1 => Si_6,                    -- added for test insertion
        out1 => Si_6_sig                -- added for test insertion
    );                                  -- added for test insertion
pout_6515: ENTITY WORK.pout             -- added for test insertion
    PORT MAP (                          -- added for test insertion
        in1 => So_1_sig,                -- added for test insertion
        out1 => So_1                    -- added for test insertion
    );                                  -- added for test insertion
pout_6516: ENTITY WORK.pout             -- added for test insertion
    PORT MAP (                          -- added for test insertion
        in1 => So_2_sig,                -- added for test insertion
        out1 => So_2                    -- added for test insertion
    );                                  -- added for test insertion
pout_6517: ENTITY WORK.pout             -- added for test insertion
    PORT MAP (                          -- added for test insertion
        in1 => So_3_sig,                -- added for test insertion
        out1 => So_3                    -- added for test insertion
    );                                  -- added for test insertion
pout_6518: ENTITY WORK.pout             -- added for test insertion
    PORT MAP (                          -- added for test insertion
        in1 => So_4_sig,                -- added for test insertion
        out1 => So_4                    -- added for test insertion
    );                                  -- added for test insertion
END ARCHITECTURE arch;
