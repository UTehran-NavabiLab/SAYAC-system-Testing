module LGC(clk, rst, readyMEM, dataBusIn, p1TRF, p2TRF, readMM, writeMM, dataBusOut, addrBus, outMuxrs1, outMuxrs2, outMuxrd, inDataTRF, writeTRF, readInst);

wire S0;
wire S1;
wire S2;
wire S3;
wire S4;
wire S5;
wire S6;
wire S7;
wire S8;
wire S9;
wire S10;
wire S11;
wire S12;
wire S13;
wire S14;
wire S15;
wire S16;
wire S17;
wire S18;
wire S19;
wire S20;
wire S21;
wire S22;
wire S23;
wire S24;
wire S25;
wire S26;
wire S27;
wire S28;
wire S29;
wire S30;
wire S31;
wire S32;
wire S33;
wire S34;
wire S35;
wire S36;
wire S37;
wire S38;
wire S39;
wire S40;
wire S41;
wire S42;
wire S43;
wire S44;
wire S45;
wire S46;
wire S47;
wire S48;
wire S49;
wire S50;
wire S51;
wire S52;
wire S53;
wire S54;
wire S55;
wire S56;
wire S57;
wire S58;
wire S59;
wire S60;
wire S61;
wire S62;
wire S63;
wire S64;
wire S65;
wire S66;
wire S67;
wire S68;
wire S69;
wire S70;
wire S71;
wire S72;
wire S73;
wire S74;
wire S75;
wire S76;
wire S77;
wire S78;
wire S79;
wire S80;
wire S81;
wire S82;
wire S83;
wire S84;
wire S85;
wire S86;
wire S87;
wire S88;
wire S89;
wire S90;
wire S91;
wire S92;
wire S93;
wire S94;
wire S95;
wire S96;
wire S97;
wire S98;
wire S99;
wire S100;
wire S101;
wire S102;
wire S103;
wire S104;
wire S105;
wire S106;
wire S107;
wire S108;
wire S109;
wire S110;
wire S111;
wire S112;
wire S113;
wire S114;
wire S115;
wire S116;
wire S117;
wire S118;
wire S119;
wire S120;
wire S121;
wire S122;
wire S123;
wire S124;
wire S125;
wire S126;
wire S127;
wire S128;
wire S129;
wire S130;
wire S131;
wire S132;
wire S133;
wire S134;
wire S135;
wire S136;
wire S137;
wire S138;
wire S139;
wire S140;
wire S141;
wire S142;
wire S143;
wire S144;
wire S145;
wire S146;
wire S147;
wire S148;
wire S149;
wire S150;
wire S151;
wire S152;
wire S153;
wire S154;
wire S155;
wire S156;
wire S157;
wire S158;
wire S159;
wire S160;
wire S161;
wire S162;
wire S163;
wire S164;
wire S165;
wire S166;
wire S167;
wire S168;
wire S169;
wire S170;
wire S171;
wire S172;
wire S173;
wire S174;
wire S175;
wire S176;
wire S177;
wire S178;
wire S179;
wire S180;
wire S181;
wire S182;
wire S183;
wire S184;
wire S185;
wire S186;
wire S187;
wire S188;
wire S189;
wire S190;
wire S191;
wire S192;
wire S193;
wire S194;
wire S195;
wire S196;
wire S197;
wire S198;
wire S199;
wire S200;
wire S201;
wire S202;
wire S203;
wire S204;
wire S205;
wire S206;
wire S207;
wire S208;
wire S209;
wire S210;
wire S211;
wire S212;
wire S213;
wire S214;
wire S215;
wire S216;
wire S217;
wire S218;
wire S219;
wire S220;
wire S221;
wire S222;
wire S223;
wire S224;
wire S225;
wire S226;
wire S227;
wire S228;
wire S229;
wire S230;
wire S231;
wire S232;
wire S233;
wire S234;
wire S235;
wire S236;
wire S237;
wire S238;
wire S239;
wire S240;
wire S241;
wire S242;
wire S243;
wire S244;
wire S245;
wire S246;
wire S247;
wire S248;
wire S249;
wire S250;
wire S251;
wire S252;
wire S253;
wire S254;
wire S255;
wire S256;
wire S257;
wire S258;
wire S259;
wire S260;
wire S261;
wire S262;
wire S263;
wire S264;
wire S265;
wire S266;
wire S267;
wire S268;
wire S269;
wire S270;
wire S271;
wire S272;
wire S273;
wire S274;
wire S275;
wire S276;
wire S277;
wire S278;
wire S279;
wire S280;
wire S281;
wire S282;
wire S283;
wire S284;
wire S285;
wire S286;
wire S287;
wire S288;
wire S289;
wire S290;
wire S291;
wire S292;
wire S293;
wire S294;
wire S295;
wire S296;
wire S297;
wire S298;
wire S299;
wire S300;
wire S301;
wire S302;
wire S303;
wire S304;
wire S305;
wire S306;
wire S307;
wire S308;
wire S309;
wire S310;
wire S311;
wire S312;
wire S313;
wire S314;
wire S315;
wire S316;
wire S317;
wire S318;
wire S319;
wire S320;
wire S321;
wire S322;
wire S323;
wire S324;
wire S325;
wire S326;
wire S327;
wire S328;
wire S329;
wire S330;
wire S331;
wire S332;
wire S333;
wire S334;
wire S335;
wire S336;
wire S337;
wire S338;
wire S339;
wire S340;
wire S341;
wire S342;
wire S343;
wire S344;
wire S345;
wire S346;
wire S347;
wire S348;
wire S349;
wire S350;
wire S351;
wire S352;
wire S353;
wire S354;
wire S355;
wire S356;
wire S357;
wire S358;
wire S359;
wire S360;
wire S361;
wire S362;
wire S363;
wire S364;
wire S365;
wire S366;
wire S367;
wire S368;
wire S369;
wire S370;
wire S371;
wire S372;
wire S373;
wire S374;
wire S375;
wire S376;
wire S377;
wire S378;
wire S379;
wire S380;
wire S381;
wire S382;
wire S383;
wire S384;
wire S385;
wire S386;
wire S387;
wire S388;
wire S389;
wire S390;
wire S391;
wire S392;
wire S393;
wire S394;
wire S395;
wire S396;
wire S397;
wire S398;
wire S399;
wire S400;
wire S401;
wire S402;
wire S403;
wire S404;
wire S405;
wire S406;
wire S407;
wire S408;
wire S409;
wire S410;
wire S411;
wire S412;
wire S413;
wire S414;
wire S415;
wire S416;
wire S417;
wire S418;
wire S419;
wire S420;
wire S421;
wire S422;
wire S423;
wire S424;
wire S425;
wire S426;
wire S427;
wire S428;
wire S429;
wire S430;
wire S431;
wire S432;
wire S433;
wire S434;
wire S435;
wire S436;
wire S437;
wire S438;
wire S439;
wire S440;
wire S441;
wire S442;
wire S443;
wire S444;
wire S445;
wire S446;
wire S447;
wire S448;
wire S449;
wire S450;
wire S451;
wire S452;
wire S453;
wire S454;
wire S455;
wire S456;
wire S457;
wire S458;
wire S459;
wire S460;
wire S461;
wire S462;
wire S463;
wire S464;
wire S465;
wire S466;
wire S467;
wire S468;
wire S469;
wire S470;
wire S471;
wire S472;
wire S473;
wire S474;
wire S475;
wire S476;
wire S477;
wire S478;
wire S479;
wire S480;
wire S481;
wire S482;
wire S483;
wire S484;
wire S485;
wire S486;
wire S487;
wire S488;
wire S489;
wire S490;
wire S491;
wire S492;
wire S493;
wire S494;
wire S495;
wire S496;
wire S497;
wire S498;
wire S499;
wire S500;
wire S501;
wire S502;
wire S503;
wire S504;
wire S505;
wire S506;
wire S507;
wire S508;
wire S509;
wire S510;
wire S511;
wire S512;
wire S513;
wire S514;
wire S515;
wire S516;
wire S517;
wire S518;
wire S519;
wire S520;
wire S521;
wire S522;
wire S523;
wire S524;
wire S525;
wire S526;
wire S527;
wire S528;
wire S529;
wire S530;
wire S531;
wire S532;
wire S533;
wire S534;
wire S535;
wire S536;
wire S537;
wire S538;
wire S539;
wire S540;
wire S541;
wire S542;
wire S543;
wire S544;
wire S545;
wire S546;
wire S547;
wire S548;
wire S549;
wire S550;
wire S551;
wire S552;
wire S553;
wire S554;
wire S555;
wire S556;
wire S557;
wire S558;
wire S559;
wire S560;
wire S561;
wire S562;
wire S563;
wire S564;
wire S565;
wire S566;
wire S567;
wire S568;
wire S569;
wire S570;
wire S571;
wire S572;
wire S573;
wire S574;
wire S575;
wire S576;
wire S577;
wire S578;
wire S579;
wire S580;
wire S581;
wire S582;
wire S583;
wire S584;
wire S585;
wire S586;
wire S587;
wire S588;
wire S589;
wire S590;
wire S591;
wire S592;
wire S593;
wire S594;
wire S595;
wire S596;
wire S597;
wire S598;
wire S599;
wire S600;
wire S601;
wire S602;
wire S603;
wire S604;
wire S605;
wire S606;
wire S607;
wire S608;
wire S609;
wire S610;
wire S611;
wire S612;
wire S613;
wire S614;
wire S615;
wire S616;
wire S617;
wire S618;
wire S619;
wire S620;
wire S621;
wire S622;
wire S623;
wire S624;
wire S625;
wire S626;
wire S627;
wire S628;
wire S629;
wire S630;
wire S631;
wire S632;
wire S633;
wire S634;
wire S635;
wire S636;
wire S637;
wire S638;
wire S639;
wire S640;
wire S641;
wire S642;
wire S643;
wire S644;
wire S645;
wire S646;
wire S647;
wire S648;
wire S649;
wire S650;
wire S651;
wire S652;
wire S653;
wire S654;
wire S655;
wire S656;
wire S657;
wire S658;
wire S659;
wire S660;
wire S661;
wire S662;
wire S663;
wire S664;
wire S665;
wire S666;
wire S667;
wire S668;
wire S669;
wire S670;
wire S671;
wire S672;
wire S673;
wire S674;
wire S675;
wire S676;
wire S677;
wire S678;
wire S679;
wire S680;
wire S681;
wire S682;
wire S683;
wire S684;
wire S685;
wire S686;
wire S687;
wire S688;
wire S689;
wire S690;
wire S691;
wire S692;
wire S693;
wire S694;
wire S695;
wire S696;
wire S697;
wire S698;
wire S699;
wire S700;
wire S701;
wire S702;
wire S703;
wire S704;
wire S705;
wire S706;
wire S707;
wire S708;
wire S709;
wire S710;
wire S711;
wire S712;
wire S713;
wire S714;
wire S715;
wire S716;
wire S717;
wire S718;
wire S719;
wire S720;
wire S721;
wire S722;
wire S723;
wire S724;
wire S725;
wire S726;
wire S727;
wire S728;
wire S729;
wire S730;
wire S731;
wire S732;
wire S733;
wire S734;
wire S735;
wire S736;
wire S737;
wire S738;
wire S739;
wire S740;
wire S741;
wire S742;
wire S743;
wire S744;
wire S745;
wire S746;
wire S747;
wire S748;
wire S749;
wire S750;
wire S751;
wire S752;
wire S753;
wire S754;
wire S755;
wire S756;
wire S757;
wire S758;
wire S759;
wire S760;
wire S761;
wire S762;
wire S763;
wire S764;
wire S765;
wire S766;
wire S767;
wire S768;
wire S769;
wire S770;
wire S771;
wire S772;
wire S773;
wire S774;
wire S775;
wire S776;
wire S777;
wire S778;
wire S779;
wire S780;
wire S781;
wire S782;
wire S783;
wire S784;
wire S785;
wire S786;
wire S787;
wire S788;
wire S789;
wire S790;
wire S791;
wire S792;
wire S793;
wire S794;
wire S795;
wire S796;
wire S797;
wire S798;
wire S799;
wire S800;
wire S801;
wire S802;
wire S803;
wire S804;
wire S805;
wire S806;
wire S807;
wire S808;
wire S809;
wire S810;
wire S811;
wire S812;
wire S813;
wire S814;
wire S815;
wire S816;
wire S817;
wire S818;
wire S819;
wire S820;
wire S821;
wire S822;
wire S823;
wire S824;
wire S825;
wire S826;
wire S827;
wire S828;
wire S829;
wire S830;
wire S831;
wire S832;
wire S833;
wire S834;
wire S835;
wire S836;
wire S837;
wire S838;
wire S839;
wire S840;
wire S841;
wire S842;
wire S843;
wire S844;
wire S845;
wire S846;
wire S847;
wire S848;
wire S849;
wire S850;
wire S851;
wire S852;
wire S853;
wire S854;
wire S855;
wire S856;
wire S857;
wire S858;
wire S859;
wire S860;
wire S861;
wire S862;
wire S863;
wire S864;
wire S865;
wire S866;
wire S867;
wire S868;
wire S869;
wire S870;
wire S871;
wire S872;
wire S873;
wire S874;
wire S875;
wire S876;
wire S877;
wire S878;
wire S879;
wire S880;
wire S881;
wire S882;
wire S883;
wire S884;
wire S885;
wire S886;
wire S887;
wire S888;
wire S889;
wire S890;
wire S891;
wire S892;
wire S893;
wire S894;
wire S895;
wire S896;
wire S897;
wire S898;
wire S899;
wire S900;
wire S901;
wire S902;
wire S903;
wire S904;
wire S905;
wire S906;
wire S907;
wire S908;
wire S909;
wire S910;
wire S911;
wire S912;
wire S913;
wire S914;
wire S915;
wire S916;
wire S917;
wire S918;
wire S919;
wire S920;
wire S921;
wire S922;
wire S923;
wire S924;
wire S925;
wire S926;
wire S927;
wire S928;
wire S929;
wire S930;
wire S931;
wire S932;
wire S933;
wire S934;
wire S935;
wire S936;
wire S937;
wire S938;
wire S939;
wire S940;
wire S941;
wire S942;
wire S943;
wire S944;
wire S945;
wire S946;
wire S947;
wire S948;
wire S949;
wire S950;
wire S951;
wire S952;
wire S953;
wire S954;
wire S955;
wire S956;
wire S957;
wire S958;
wire S959;
wire S960;
wire S961;
wire S962;
wire S963;
wire S964;
wire S965;
wire S966;
wire S967;
wire S968;
wire S969;
wire S970;
wire S971;
wire S972;
wire S973;
wire S974;
wire S975;
wire S976;
wire S977;
wire S978;
wire S979;
wire S980;
wire S981;
wire S982;
wire S983;
wire S984;
wire S985;
wire S986;
wire S987;
wire S988;
wire S989;
wire S990;
wire S991;
wire S992;
wire S993;
wire S994;
wire S995;
wire S996;
wire S997;
wire S998;
wire S999;
wire S1000;
wire S1001;
wire S1002;
wire S1003;
wire S1004;
wire S1005;
wire S1006;
wire S1007;
wire S1008;
wire S1009;
wire S1010;
wire S1011;
wire S1012;
wire S1013;
wire S1014;
wire S1015;
wire S1016;
wire S1017;
wire S1018;
wire S1019;
wire S1020;
wire S1021;
wire S1022;
wire S1023;
wire S1024;
wire S1025;
wire S1026;
wire S1027;
wire S1028;
wire S1029;
wire S1030;
wire S1031;
wire S1032;
wire S1033;
wire S1034;
wire S1035;
wire S1036;
wire S1037;
wire S1038;
wire S1039;
wire S1040;
wire S1041;
wire S1042;
wire S1043;
wire S1044;
wire S1045;
wire S1046;
wire S1047;
wire S1048;
wire S1049;
wire S1050;
wire S1051;
wire S1052;
wire S1053;
wire S1054;
wire S1055;
wire S1056;
wire S1057;
wire S1058;
wire S1059;
wire S1060;
wire S1061;
wire S1062;
wire S1063;
wire S1064;
wire S1065;
wire S1066;
wire S1067;
wire S1068;
wire S1069;
wire S1070;
wire S1071;
wire S1072;
wire S1073;
wire S1074;
wire S1075;
wire S1076;
wire S1077;
wire S1078;
wire S1079;
wire S1080;
wire S1081;
wire S1082;
wire S1083;
wire S1084;
wire S1085;
wire S1086;
wire S1087;
wire S1088;
wire S1089;
wire S1090;
wire S1091;
wire S1092;
wire S1093;
wire S1094;
wire S1095;
wire S1096;
wire S1097;
wire S1098;
wire S1099;
wire S1100;
wire S1101;
wire S1102;
wire S1103;
wire S1104;
wire S1105;
wire S1106;
wire S1107;
wire S1108;
wire S1109;
wire S1110;
wire S1111;
wire S1112;
wire S1113;
wire S1114;
wire S1115;
wire S1116;
wire S1117;
wire S1118;
wire S1119;
wire S1120;
wire S1121;
wire S1122;
wire S1123;
wire S1124;
wire S1125;
wire S1126;
wire S1127;
wire S1128;
wire S1129;
wire S1130;
wire S1131;
wire S1132;
wire S1133;
wire S1134;
wire S1135;
wire S1136;
wire S1137;
wire S1138;
wire S1139;
wire S1140;
wire S1141;
wire S1142;
wire S1143;
wire S1144;
wire S1145;
wire S1146;
wire S1147;
wire S1148;
wire S1149;
wire S1150;
wire S1151;
wire S1152;
wire S1153;
wire S1154;
wire S1155;
wire S1156;
wire S1157;
wire S1158;
wire S1159;
wire S1160;
wire S1161;
wire S1162;
wire S1163;
wire S1164;
wire S1165;
wire S1166;
wire S1167;
wire S1168;
wire S1169;
wire S1170;
wire S1171;
wire S1172;
wire S1173;
wire S1174;
wire S1175;
wire S1176;
wire S1177;
wire S1178;
wire S1179;
wire S1180;
wire S1181;
wire S1182;
wire S1183;
wire S1184;
wire S1185;
wire S1186;
wire S1187;
wire S1188;
wire S1189;
wire S1190;
wire S1191;
wire S1192;
wire S1193;
wire S1194;
wire S1195;
wire S1196;
wire S1197;
wire S1198;
wire S1199;
wire S1200;
wire S1201;
wire S1202;
wire S1203;
wire S1204;
wire S1205;
wire S1206;
wire S1207;
wire S1208;
wire S1209;
wire S1210;
wire S1211;
wire S1212;
wire S1213;
wire S1214;
wire S1215;
wire S1216;
wire S1217;
wire S1218;
wire S1219;
wire S1220;
wire S1221;
wire S1222;
wire S1223;
wire S1224;
wire S1225;
wire S1226;
wire S1227;
wire S1228;
wire S1229;
wire S1230;
wire S1231;
wire S1232;
wire S1233;
wire S1234;
wire S1235;
wire S1236;
wire S1237;
wire S1238;
wire S1239;
wire S1240;
wire S1241;
wire S1242;
wire S1243;
wire S1244;
wire S1245;
wire S1246;
wire S1247;
wire S1248;
wire S1249;
wire S1250;
wire S1251;
wire S1252;
wire S1253;
wire S1254;
wire S1255;
wire S1256;
wire S1257;
wire S1258;
wire S1259;
wire S1260;
wire S1261;
wire S1262;
wire S1263;
wire S1264;
wire S1265;
wire S1266;
wire S1267;
wire S1268;
wire S1269;
wire S1270;
wire S1271;
wire S1272;
wire S1273;
wire S1274;
wire S1275;
wire S1276;
wire S1277;
wire S1278;
wire S1279;
wire S1280;
wire S1281;
wire S1282;
wire S1283;
wire S1284;
wire S1285;
wire S1286;
wire S1287;
wire S1288;
wire S1289;
wire S1290;
wire S1291;
wire S1292;
wire S1293;
wire S1294;
wire S1295;
wire S1296;
wire S1297;
wire S1298;
wire S1299;
wire S1300;
wire S1301;
wire S1302;
wire S1303;
wire S1304;
wire S1305;
wire S1306;
wire S1307;
wire S1308;
wire S1309;
wire S1310;
wire S1311;
wire S1312;
wire S1313;
wire S1314;
wire S1315;
wire S1316;
wire S1317;
wire S1318;
wire S1319;
wire S1320;
wire S1321;
wire S1322;
wire S1323;
wire S1324;
wire S1325;
wire S1326;
wire S1327;
wire S1328;
wire S1329;
wire S1330;
wire S1331;
wire S1332;
wire S1333;
wire S1334;
wire S1335;
wire S1336;
wire S1337;
wire S1338;
wire S1339;
wire S1340;
wire S1341;
wire S1342;
wire S1343;
wire S1344;
wire S1345;
wire S1346;
wire S1347;
wire S1348;
wire S1349;
wire S1350;
wire S1351;
wire S1352;
wire S1353;
wire S1354;
wire S1355;
wire S1356;
wire S1357;
wire S1358;
wire S1359;
wire S1360;
wire S1361;
wire S1362;
wire S1363;
wire S1364;
wire S1365;
wire S1366;
wire S1367;
wire S1368;
wire S1369;
wire S1370;
wire S1371;
wire S1372;
wire S1373;
wire S1374;
wire S1375;
wire S1376;
wire S1377;
wire S1378;
wire S1379;
wire S1380;
wire S1381;
wire S1382;
wire S1383;
wire S1384;
wire S1385;
wire S1386;
wire S1387;
wire S1388;
wire S1389;
wire S1390;
wire S1391;
wire S1392;
wire S1393;
wire S1394;
wire S1395;
wire S1396;
wire S1397;
wire S1398;
wire S1399;
wire S1400;
wire S1401;
wire S1402;
wire S1403;
wire S1404;
wire S1405;
wire S1406;
wire S1407;
wire S1408;
wire S1409;
wire S1410;
wire S1411;
wire S1412;
wire S1413;
wire S1414;
wire S1415;
wire S1416;
wire S1417;
wire S1418;
wire S1419;
wire S1420;
wire S1421;
wire S1422;
wire S1423;
wire S1424;
wire S1425;
wire S1426;
wire S1427;
wire S1428;
wire S1429;
wire S1430;
wire S1431;
wire S1432;
wire S1433;
wire S1434;
wire S1435;
wire S1436;
wire S1437;
wire S1438;
wire S1439;
wire S1440;
wire S1441;
wire S1442;
wire S1443;
wire S1444;
wire S1445;
wire S1446;
wire S1447;
wire S1448;
wire S1449;
wire S1450;
wire S1451;
wire S1452;
wire S1453;
wire S1454;
wire S1455;
wire S1456;
wire S1457;
wire S1458;
wire S1459;
wire S1460;
wire S1461;
wire S1462;
wire S1463;
wire S1464;
wire S1465;
wire S1466;
wire S1467;
wire S1468;
wire S1469;
wire S1470;
wire S1471;
wire S1472;
wire S1473;
wire S1474;
wire S1475;
wire S1476;
wire S1477;
wire S1478;
wire S1479;
wire S1480;
wire S1481;
wire S1482;
wire S1483;
wire S1484;
wire S1485;
wire S1486;
wire S1487;
wire S1488;
wire S1489;
wire S1490;
wire S1491;
wire S1492;
wire S1493;
wire S1494;
wire S1495;
wire S1496;
wire S1497;
wire S1498;
wire S1499;
wire S1500;
wire S1501;
wire S1502;
wire S1503;
wire S1504;
wire S1505;
wire S1506;
wire S1507;
wire S1508;
wire S1509;
wire S1510;
wire S1511;
wire S1512;
wire S1513;
wire S1514;
wire S1515;
wire S1516;
wire S1517;
wire S1518;
wire S1519;
wire S1520;
wire S1521;
wire S1522;
wire S1523;
wire S1524;
wire S1525;
wire S1526;
wire S1527;
wire S1528;
wire S1529;
wire S1530;
wire S1531;
wire S1532;
wire S1533;
wire S1534;
wire S1535;
wire S1536;
wire S1537;
wire S1538;
wire S1539;
wire S1540;
wire S1541;
wire S1542;
wire S1543;
wire S1544;
wire S1545;
wire S1546;
wire S1547;
wire S1548;
wire S1549;
wire S1550;
wire S1551;
wire S1552;
wire S1553;
wire S1554;
wire S1555;
wire S1556;
wire S1557;
wire S1558;
wire S1559;
wire S1560;
wire S1561;
wire S1562;
wire S1563;
wire S1564;
wire S1565;
wire S1566;
wire S1567;
wire S1568;
wire S1569;
wire S1570;
wire S1571;
wire S1572;
wire S1573;
wire S1574;
wire S1575;
wire S1576;
wire S1577;
wire S1578;
wire S1579;
wire S1580;
wire S1581;
wire S1582;
wire S1583;
wire S1584;
wire S1585;
wire S1586;
wire S1587;
wire S1588;
wire S1589;
wire S1590;
wire S1591;
wire S1592;
wire S1593;
wire S1594;
wire S1595;
wire S1596;
wire S1597;
wire S1598;
wire S1599;
wire S1600;
wire S1601;
wire S1602;
wire S1603;
wire S1604;
wire S1605;
wire S1606;
wire S1607;
wire S1608;
wire S1609;
wire S1610;
wire S1611;
wire S1612;
wire S1613;
wire S1614;
wire S1615;
wire S1616;
wire S1617;
wire S1618;
wire S1619;
wire S1620;
wire S1621;
wire S1622;
wire S1623;
wire S1624;
wire S1625;
wire S1626;
wire S1627;
wire S1628;
wire S1629;
wire S1630;
wire S1631;
wire S1632;
wire S1633;
wire S1634;
wire S1635;
wire S1636;
wire S1637;
wire S1638;
wire S1639;
wire S1640;
wire S1641;
wire S1642;
wire S1643;
wire S1644;
wire S1645;
wire S1646;
wire S1647;
wire S1648;
wire S1649;
wire S1650;
wire S1651;
wire S1652;
wire S1653;
wire S1654;
wire S1655;
wire S1656;
wire S1657;
wire S1658;
wire S1659;
wire S1660;
wire S1661;
wire S1662;
wire S1663;
wire S1664;
wire S1665;
wire S1666;
wire S1667;
wire S1668;
wire S1669;
wire S1670;
wire S1671;
wire S1672;
wire S1673;
wire S1674;
wire S1675;
wire S1676;
wire S1677;
wire S1678;
wire S1679;
wire S1680;
wire S1681;
wire S1682;
wire S1683;
wire S1684;
wire S1685;
wire S1686;
wire S1687;
wire S1688;
wire S1689;
wire S1690;
wire S1691;
wire S1692;
wire S1693;
wire S1694;
wire S1695;
wire S1696;
wire S1697;
wire S1698;
wire S1699;
wire S1700;
wire S1701;
wire S1702;
wire S1703;
wire S1704;
wire S1705;
wire S1706;
wire S1707;
wire S1708;
wire S1709;
wire S1710;
wire S1711;
wire S1712;
wire S1713;
wire S1714;
wire S1715;
wire S1716;
wire S1717;
wire S1718;
wire S1719;
wire S1720;
wire S1721;
wire S1722;
wire S1723;
wire S1724;
wire S1725;
wire S1726;
wire S1727;
wire S1728;
wire S1729;
wire S1730;
wire S1731;
wire S1732;
wire S1733;
wire S1734;
wire S1735;
wire S1736;
wire S1737;
wire S1738;
wire S1739;
wire S1740;
wire S1741;
wire S1742;
wire S1743;
wire S1744;
wire S1745;
wire S1746;
wire S1747;
wire S1748;
wire S1749;
wire S1750;
wire S1751;
wire S1752;
wire S1753;
wire S1754;
wire S1755;
wire S1756;
wire S1757;
wire S1758;
wire S1759;
wire S1760;
wire S1761;
wire S1762;
wire S1763;
wire S1764;
wire S1765;
wire S1766;
wire S1767;
wire S1768;
wire S1769;
wire S1770;
wire S1771;
wire S1772;
wire S1773;
wire S1774;
wire S1775;
wire S1776;
wire S1777;
wire S1778;
wire S1779;
wire S1780;
wire S1781;
wire S1782;
wire S1783;
wire S1784;
wire S1785;
wire S1786;
wire S1787;
wire S1788;
wire S1789;
wire S1790;
wire S1791;
wire S1792;
wire S1793;
wire S1794;
wire S1795;
wire S1796;
wire S1797;
wire S1798;
wire S1799;
wire S1800;
wire S1801;
wire S1802;
wire S1803;
wire S1804;
wire S1805;
wire S1806;
wire S1807;
wire S1808;
wire S1809;
wire S1810;
wire S1811;
wire S1812;
wire S1813;
wire S1814;
wire S1815;
wire S1816;
wire S1817;
wire S1818;
wire S1819;
wire S1820;
wire S1821;
wire S1822;
wire S1823;
wire S1824;
wire S1825;
wire S1826;
wire S1827;
wire S1828;
wire S1829;
wire S1830;
wire S1831;
wire S1832;
wire S1833;
wire S1834;
wire S1835;
wire S1836;
wire S1837;
wire S1838;
wire S1839;
wire S1840;
wire S1841;
wire S1842;
wire S1843;
wire S1844;
wire S1845;
wire S1846;
wire S1847;
wire S1848;
wire S1849;
wire S1850;
wire S1851;
wire S1852;
wire S1853;
wire S1854;
wire S1855;
wire S1856;
wire S1857;
wire S1858;
wire S1859;
wire S1860;
wire S1861;
wire S1862;
wire S1863;
wire S1864;
wire S1865;
wire S1866;
wire S1867;
wire S1868;
wire S1869;
wire S1870;
wire S1871;
wire S1872;
wire S1873;
wire S1874;
wire S1875;
wire S1876;
wire S1877;
wire S1878;
wire S1879;
wire S1880;
wire S1881;
wire S1882;
wire S1883;
wire S1884;
wire S1885;
wire S1886;
wire S1887;
wire S1888;
wire S1889;
wire S1890;
wire S1891;
wire S1892;
wire S1893;
wire S1894;
wire S1895;
wire S1896;
wire S1897;
wire S1898;
wire S1899;
wire S1900;
wire S1901;
wire S1902;
wire S1903;
wire S1904;
wire S1905;
wire S1906;
wire S1907;
wire S1908;
wire S1909;
wire S1910;
wire S1911;
wire S1912;
wire S1913;
wire S1914;
wire S1915;
wire S1916;
wire S1917;
wire S1918;
wire S1919;
wire S1920;
wire S1921;
wire S1922;
wire S1923;
wire S1924;
wire S1925;
wire S1926;
wire S1927;
wire S1928;
wire S1929;
wire S1930;
wire S1931;
wire S1932;
wire S1933;
wire S1934;
wire S1935;
wire S1936;
wire S1937;
wire S1938;
wire S1939;
wire S1940;
wire S1941;
wire S1942;
wire S1943;
wire S1944;
wire S1945;
wire S1946;
wire S1947;
wire S1948;
wire S1949;
wire S1950;
wire S1951;
wire S1952;
wire S1953;
wire S1954;
wire S1955;
wire S1956;
wire S1957;
wire S1958;
wire S1959;
wire S1960;
wire S1961;
wire S1962;
wire S1963;
wire S1964;
wire S1965;
wire S1966;
wire S1967;
wire S1968;
wire S1969;
wire S1970;
wire S1971;
wire S1972;
wire S1973;
wire S1974;
wire S1975;
wire S1976;
wire S1977;
wire S1978;
wire S1979;
wire S1980;
wire S1981;
wire S1982;
wire S1983;
wire S1984;
wire S1985;
wire S1986;
wire S1987;
wire S1988;
wire S1989;
wire S1990;
wire S1991;
wire S1992;
wire S1993;
wire S1994;
wire S1995;
wire S1996;
wire S1997;
wire S1998;
wire S1999;
wire S2000;
wire S2001;
wire S2002;
wire S2003;
wire S2004;
wire S2005;
wire S2006;
wire S2007;
wire S2008;
wire S2009;
wire S2010;
wire S2011;
wire S2012;
wire S2013;
wire S2014;
wire S2015;
wire S2016;
wire S2017;
wire S2018;
wire S2019;
wire S2020;
wire S2021;
wire S2022;
wire S2023;
wire S2024;
wire S2025;
wire S2026;
wire S2027;
wire S2028;
wire S2029;
wire S2030;
wire S2031;
wire S2032;
wire S2033;
wire S2034;
wire S2035;
wire S2036;
wire S2037;
wire S2038;
wire S2039;
wire S2040;
wire S2041;
wire S2042;
wire S2043;
wire S2044;
wire S2045;
wire S2046;
wire S2047;
wire S2048;
wire S2049;
wire S2050;
wire S2051;
wire S2052;
wire S2053;
wire S2054;
wire S2055;
wire S2056;
wire S2057;
wire S2058;
wire S2059;
wire S2060;
wire S2061;
wire S2062;
wire S2063;
wire S2064;
wire S2065;
wire S2066;
wire S2067;
wire S2068;
wire S2069;
wire S2070;
wire S2071;
wire S2072;
wire S2073;
wire S2074;
wire S2075;
wire S2076;
wire S2077;
wire S2078;
wire S2079;
wire S2080;
wire S2081;
wire S2082;
wire S2083;
wire S2084;
wire S2085;
wire S2086;
wire S2087;
wire S2088;
wire S2089;
wire S2090;
wire S2091;
wire S2092;
wire S2093;
wire S2094;
wire S2095;
wire S2096;
wire S2097;
wire S2098;
wire S2099;
wire S2100;
wire S2101;
wire S2102;
wire S2103;
wire S2104;
wire S2105;
wire S2106;
wire S2107;
wire S2108;
wire S2109;
wire S2110;
wire S2111;
wire S2112;
wire S2113;
wire S2114;
wire S2115;
wire S2116;
wire S2117;
wire S2118;
wire S2119;
wire S2120;
wire S2121;
wire S2122;
wire S2123;
wire S2124;
wire S2125;
wire S2126;
wire S2127;
wire S2128;
wire S2129;
wire S2130;
wire S2131;
wire S2132;
wire S2133;
wire S2134;
wire S2135;
wire S2136;
wire S2137;
wire S2138;
wire S2139;
wire S2140;
wire S2141;
wire S2142;
wire S2143;
wire S2144;
wire S2145;
wire S2146;
wire S2147;
wire S2148;
wire S2149;
wire S2150;
wire S2151;
wire S2152;
wire S2153;
wire S2154;
wire S2155;
wire S2156;
wire S2157;
wire S2158;
wire S2159;
wire S2160;
wire S2161;
wire S2162;
wire S2163;
wire S2164;
wire S2165;
wire S2166;
wire S2167;
wire S2168;
wire S2169;
wire S2170;
wire S2171;
wire S2172;
wire S2173;
wire S2174;
wire S2175;
wire S2176;
wire S2177;
wire S2178;
wire S2179;
wire S2180;
wire S2181;
wire S2182;
wire S2183;
wire S2184;
wire S2185;
wire S2186;
wire S2187;
wire S2188;
wire S2189;
wire S2190;
wire S2191;
wire S2192;
wire S2193;
wire S2194;
wire S2195;
wire S2196;
wire S2197;
wire S2198;
wire S2199;
wire S2200;
wire S2201;
wire S2202;
wire S2203;
wire S2204;
wire S2205;
wire S2206;
wire S2207;
wire S2208;
wire S2209;
wire S2210;
wire S2211;
wire S2212;
wire S2213;
wire S2214;
wire S2215;
wire S2216;
wire S2217;
wire S2218;
wire S2219;
wire S2220;
wire S2221;
wire S2222;
wire S2223;
wire S2224;
wire S2225;
wire S2226;
wire S2227;
wire S2228;
wire S2229;
wire S2230;
wire S2231;
wire S2232;
wire S2233;
wire S2234;
wire S2235;
wire S2236;
wire S2237;
wire S2238;
wire S2239;
wire S2240;
wire S2241;
wire S2242;
wire S2243;
wire S2244;
wire S2245;
wire S2246;
wire S2247;
wire S2248;
wire S2249;
wire S2250;
wire S2251;
wire S2252;
wire S2253;
wire S2254;
wire S2255;
wire S2256;
wire S2257;
wire S2258;
wire S2259;
wire S2260;
wire S2261;
wire S2262;
wire S2263;
wire S2264;
wire S2265;
wire S2266;
wire S2267;
wire S2268;
wire S2269;
wire S2270;
wire S2271;
wire S2272;
wire S2273;
wire S2274;
wire S2275;
wire S2276;
wire S2277;
wire S2278;
wire S2279;
wire S2280;
wire S2281;
wire S2282;
wire S2283;
wire S2284;
wire S2285;
wire S2286;
wire S2287;
wire S2288;
wire S2289;
wire S2290;
wire S2291;
wire S2292;
wire S2293;
wire S2294;
wire S2295;
wire S2296;
wire S2297;
wire S2298;
wire S2299;
wire S2300;
wire S2301;
wire S2302;
wire S2303;
wire S2304;
wire S2305;
wire S2306;
wire S2307;
wire S2308;
wire S2309;
wire S2310;
wire S2311;
wire S2312;
wire S2313;
wire S2314;
wire S2315;
wire S2316;
wire S2317;
wire S2318;
wire S2319;
wire S2320;
wire S2321;
wire S2322;
wire S2323;
wire S2324;
wire S2325;
wire S2326;
wire S2327;
wire S2328;
wire S2329;
wire S2330;
wire S2331;
wire S2332;
wire S2333;
wire S2334;
wire S2335;
wire S2336;
wire S2337;
wire S2338;
wire S2339;
wire S2340;
wire S2341;
wire S2342;
wire S2343;
wire S2344;
wire S2345;
wire S2346;
wire S2347;
wire S2348;
wire S2349;
wire S2350;
wire S2351;
wire S2352;
wire S2353;
wire S2354;
wire S2355;
wire S2356;
wire S2357;
wire S2358;
wire S2359;
wire S2360;
wire S2361;
wire S2362;
wire S2363;
wire S2364;
wire S2365;
wire S2366;
wire S2367;
wire S2368;
wire S2369;
wire S2370;
wire S2371;
wire S2372;
wire S2373;
wire S2374;
wire S2375;
wire S2376;
wire S2377;
wire S2378;
wire S2379;
wire S2380;
wire S2381;
wire S2382;
wire S2383;
wire S2384;
wire S2385;
wire S2386;
wire S2387;
wire S2388;
wire S2389;
wire S2390;
wire S2391;
wire S2392;
wire S2393;
wire S2394;
wire S2395;
wire S2396;
wire S2397;
wire S2398;
wire S2399;
wire S2400;
wire S2401;
wire S2402;
wire S2403;
wire S2404;
wire S2405;
wire S2406;
wire S2407;
wire S2408;
wire S2409;
wire S2410;
wire S2411;
wire S2412;
wire S2413;
wire S2414;
wire S2415;
wire S2416;
wire S2417;
wire S2418;
wire S2419;
wire S2420;
wire S2421;
wire S2422;
wire S2423;
wire S2424;
wire S2425;
wire S2426;
wire S2427;
wire S2428;
wire S2429;
wire S2430;
wire S2431;
wire S2432;
wire S2433;
wire S2434;
wire S2435;
wire S2436;
wire S2437;
wire S2438;
wire S2439;
wire S2440;
wire S2441;
wire S2442;
wire S2443;
wire S2444;
wire S2445;
wire S2446;
wire S2447;
wire S2448;
wire S2449;
wire S2450;
wire S2451;
wire S2452;
wire S2453;
wire S2454;
wire S2455;
wire S2456;
wire S2457;
wire S2458;
wire S2459;
wire S2460;
wire S2461;
wire S2462;
wire S2463;
wire S2464;
wire S2465;
wire S2466;
wire S2467;
wire S2468;
wire S2469;
wire S2470;
wire S2471;
wire S2472;
wire S2473;
wire S2474;
wire S2475;
wire S2476;
wire S2477;
wire S2478;
wire S2479;
wire S2480;
wire S2481;
wire S2482;
wire S2483;
wire S2484;
wire S2485;
wire S2486;
wire S2487;
wire S2488;
wire S2489;
wire S2490;
wire S2491;
wire S2492;
wire S2493;
wire S2494;
wire S2495;
wire S2496;
wire S2497;
wire S2498;
wire S2499;
wire S2500;
wire S2501;
wire S2502;
wire S2503;
wire S2504;
wire S2505;
wire S2506;
wire S2507;
wire S2508;
wire S2509;
wire S2510;
wire S2511;
wire S2512;
wire S2513;
wire S2514;
wire S2515;
wire S2516;
wire S2517;
wire S2518;
wire S2519;
wire S2520;
wire S2521;
wire S2522;
wire S2523;
wire S2524;
wire S2525;
wire S2526;
wire S2527;
wire S2528;
wire S2529;
wire S2530;
wire S2531;
wire S2532;
wire S2533;
wire S2534;
wire S2535;
wire S2536;
wire S2537;
wire S2538;
wire S2539;
wire S2540;
wire S2541;
wire S2542;
wire S2543;
wire S2544;
wire S2545;
wire S2546;
wire S2547;
wire S2548;
wire S2549;
wire S2550;
wire S2551;
wire S2552;
wire S2553;
wire S2554;
wire S2555;
wire S2556;
wire S2557;
wire S2558;
wire S2559;
wire S2560;
wire S2561;
wire S2562;
wire S2563;
wire S2564;
wire S2565;
wire S2566;
wire S2567;
wire S2568;
wire S2569;
wire S2570;
wire S2571;
wire S2572;
wire S2573;
wire S2574;
wire S2575;
wire S2576;
wire S2577;
wire S2578;
wire S2579;
wire S2580;
wire S2581;
wire S2582;
wire S2583;
wire S2584;
wire S2585;
wire S2586;
wire S2587;
wire S2588;
wire S2589;
wire S2590;
wire S2591;
wire S2592;
wire S2593;
wire S2594;
wire S2595;
wire S2596;
wire S2597;
wire S2598;
wire S2599;
wire S2600;
wire S2601;
wire S2602;
wire S2603;
wire S2604;
wire S2605;
wire S2606;
wire S2607;
wire S2608;
wire S2609;
wire S2610;
wire S2611;
wire S2612;
wire S2613;
wire S2614;
wire S2615;
wire S2616;
wire S2617;
wire S2618;
wire S2619;
wire S2620;
wire S2621;
wire S2622;
wire S2623;
wire S2624;
wire S2625;
wire S2626;
wire S2627;
wire S2628;
wire S2629;
wire S2630;
wire S2631;
wire S2632;
wire S2633;
wire S2634;
wire S2635;
wire S2636;
wire S2637;
wire S2638;
wire S2639;
wire S2640;
wire S2641;
wire S2642;
wire S2643;
wire S2644;
wire S2645;
wire S2646;
wire S2647;
wire S2648;
wire S2649;
wire S2650;
wire S2651;
wire S2652;
wire S2653;
wire S2654;
wire S2655;
wire S2656;
wire S2657;
wire S2658;
wire S2659;
wire S2660;
wire S2661;
wire S2662;
wire S2663;
wire S2664;
wire S2665;
wire S2666;
wire S2667;
wire S2668;
wire S2669;
wire S2670;
wire S2671;
wire S2672;
wire S2673;
wire S2674;
wire S2675;
wire S2676;
wire S2677;
wire S2678;
wire S2679;
wire S2680;
wire S2681;
wire S2682;
wire S2683;
wire S2684;
wire S2685;
wire S2686;
wire S2687;
wire S2688;
wire S2689;
wire S2690;
wire S2691;
wire S2692;
wire S2693;
wire S2694;
wire S2695;
wire S2696;
wire S2697;
wire S2698;
wire S2699;
wire S2700;
wire S2701;
wire S2702;
wire S2703;
wire S2704;
wire S2705;
wire S2706;
wire S2707;
wire S2708;
wire S2709;
wire S2710;
wire S2711;
wire S2712;
wire S2713;
wire S2714;
wire S2715;
wire S2716;
wire S2717;
wire S2718;
wire S2719;
wire S2720;
wire S2721;
wire S2722;
wire S2723;
wire S2724;
wire S2725;
wire S2726;
wire S2727;
wire S2728;
wire S2729;
wire S2730;
wire S2731;
wire S2732;
wire S2733;
wire S2734;
wire S2735;
wire S2736;
wire S2737;
wire S2738;
wire S2739;
wire S2740;
wire S2741;
wire S2742;
wire S2743;
wire S2744;
wire S2745;
wire S2746;
wire S2747;
wire S2748;
wire S2749;
wire S2750;
wire S2751;
wire S2752;
wire S2753;
wire S2754;
wire S2755;
wire S2756;
wire S2757;
wire S2758;
wire S2759;
wire S2760;
wire S2761;
wire S2762;
wire S2763;
wire S2764;
wire S2765;
wire S2766;
wire S2767;
wire S2768;
wire S2769;
wire S2770;
wire S2771;
wire S2772;
wire S2773;
wire S2774;
wire S2775;
wire S2776;
wire S2777;
wire S2778;
wire S2779;
wire S2780;
wire S2781;
wire S2782;
wire S2783;
wire S2784;
wire S2785;
wire S2786;
wire S2787;
wire S2788;
wire S2789;
wire S2790;
wire S2791;
wire S2792;
wire S2793;
wire S2794;
wire S2795;
wire S2796;
wire S2797;
wire S2798;
wire S2799;
wire S2800;
wire S2801;
wire S2802;
wire S2803;
wire S2804;
wire S2805;
wire S2806;
wire S2807;
wire S2808;
wire S2809;
wire S2810;
wire S2811;
wire S2812;
wire S2813;
wire S2814;
wire S2815;
wire S2816;
wire S2817;
wire S2818;
wire S2819;
wire S2820;
wire S2821;
wire S2822;
wire S2823;
wire S2824;
wire S2825;
wire S2826;
wire S2827;
wire S2828;
wire S2829;
wire S2830;
wire S2831;
wire S2832;
wire S2833;
wire S2834;
wire S2835;
wire S2836;
wire S2837;
wire S2838;
wire S2839;
wire S2840;
wire S2841;
wire S2842;
wire S2843;
wire S2844;
wire S2845;
wire S2846;
wire S2847;
wire S2848;
wire S2849;
wire S2850;
wire S2851;
wire S2852;
wire S2853;
wire S2854;
wire S2855;
wire S2856;
wire S2857;
wire S2858;
wire S2859;
wire S2860;
wire S2861;
wire S2862;
wire S2863;
wire S2864;
wire S2865;
wire S2866;
wire S2867;
wire S2868;
wire S2869;
wire S2870;
wire S2871;
wire S2872;
wire S2873;
wire S2874;
wire S2875;
wire S2876;
wire S2877;
wire S2878;
wire S2879;
wire S2880;
wire S2881;
wire S2882;
wire S2883;
wire S2884;
wire S2885;
wire S2886;
wire S2887;
wire S2888;
wire S2889;
wire S2890;
wire S2891;
wire S2892;
wire S2893;
wire S2894;
wire S2895;
wire S2896;
wire S2897;
wire S2898;
wire S2899;
wire S2900;
wire S2901;
wire S2902;
wire S2903;
wire S2904;
wire S2905;
wire S2906;
wire S2907;
wire S2908;
wire S2909;
wire S2910;
wire S2911;
wire S2912;
wire S2913;
wire S2914;
wire S2915;
wire S2916;
wire S2917;
wire S2918;
wire S2919;
wire S2920;
wire S2921;
wire S2922;
wire S2923;
wire S2924;
wire S2925;
wire S2926;
wire S2927;
wire S2928;
wire S2929;
wire S2930;
wire S2931;
wire S2932;
wire S2933;
wire S2934;
wire S2935;
wire S2936;
wire S2937;
wire S2938;
wire S2939;
wire S2940;
wire S2941;
wire S2942;
wire S2943;
wire S2944;
wire S2945;
wire S2946;
wire S2947;
wire S2948;
wire S2949;
wire S2950;
wire S2951;
wire S2952;
wire S2953;
wire S2954;
wire S2955;
wire S2956;
wire S2957;
wire S2958;
wire S2959;
wire S2960;
wire S2961;
wire S2962;
wire S2963;
wire S2964;
wire S2965;
wire S2966;
wire S2967;
wire S2968;
wire S2969;
wire S2970;
wire S2971;
wire S2972;
wire S2973;
wire S2974;
wire S2975;
wire S2976;
wire S2977;
wire S2978;
wire S2979;
wire S2980;
wire S2981;
wire S2982;
wire S2983;
wire S2984;
wire S2985;
wire S2986;
wire S2987;
wire S2988;
wire S2989;
wire S2990;
wire S2991;
wire S2992;
wire S2993;
wire S2994;
wire S2995;
wire S2996;
wire S2997;
wire S2998;
wire S2999;
wire S3000;
wire S3001;
wire S3002;
wire S3003;
wire S3004;
wire S3005;
wire S3006;
wire S3007;
wire S3008;
wire S3009;
wire S3010;
wire S3011;
wire S3012;
wire S3013;
wire S3014;
wire S3015;
wire S3016;
wire S3017;
wire S3018;
wire S3019;
wire S3020;
wire S3021;
wire S3022;
wire S3023;
wire S3024;
wire S3025;
wire S3026;
wire S3027;
wire S3028;
wire S3029;
wire S3030;
wire S3031;
wire S3032;
wire S3033;
wire S3034;
wire S3035;
wire S3036;
wire S3037;
wire S3038;
wire S3039;
wire S3040;
wire S3041;
wire S3042;
wire S3043;
wire S3044;
wire S3045;
wire S3046;
wire S3047;
wire S3048;
wire S3049;
wire S3050;
wire S3051;
wire S3052;
wire S3053;
wire S3054;
wire S3055;
wire S3056;
wire S3057;
wire S3058;
wire S3059;
wire S3060;
wire S3061;
wire S3062;
wire S3063;
wire S3064;
wire S3065;
wire S3066;
wire S3067;
wire S3068;
wire S3069;
wire S3070;
wire S3071;
wire S3072;
wire S3073;
wire S3074;
wire S3075;
wire S3076;
wire S3077;
wire S3078;
wire S3079;
wire S3080;
wire S3081;
wire S3082;
wire S3083;
wire S3084;
wire S3085;
wire S3086;
wire S3087;
wire S3088;
wire S3089;
wire S3090;
wire S3091;
wire S3092;
wire S3093;
wire S3094;
wire S3095;
wire S3096;
wire S3097;
wire S3098;
wire S3099;
wire S3100;
wire S3101;
wire S3102;
wire S3103;
wire S3104;
wire S3105;
wire S3106;
wire S3107;
wire S3108;
wire S3109;
wire S3110;
wire S3111;
wire S3112;
wire S3113;
wire S3114;
wire S3115;
wire S3116;
wire S3117;
wire S3118;
wire S3119;
wire S3120;
wire S3121;
wire S3122;
wire S3123;
wire S3124;
wire S3125;
wire S3126;
wire S3127;
wire S3128;
wire S3129;
wire S3130;
wire S3131;
wire S3132;
wire S3133;
wire S3134;
wire S3135;
wire S3136;
wire S3137;
wire S3138;
wire S3139;
wire S3140;
wire S3141;
wire S3142;
wire S3143;
wire S3144;
wire S3145;
wire S3146;
wire S3147;
wire S3148;
wire S3149;
wire S3150;
wire S3151;
wire S3152;
wire S3153;
wire S3154;
wire S3155;
wire S3156;
wire S3157;
wire S3158;
wire S3159;
wire S3160;
wire S3161;
wire S3162;
wire S3163;
wire S3164;
wire S3165;
wire S3166;
wire S3167;
wire S3168;
wire S3169;
wire S3170;
wire S3171;
wire S3172;
wire S3173;
wire S3174;
wire S3175;
wire S3176;
wire S3177;
wire S3178;
wire S3179;
wire S3180;
wire S3181;
wire S3182;
wire S3183;
wire S3184;
wire S3185;
wire S3186;
wire S3187;
wire S3188;
wire S3189;
wire S3190;
wire S3191;
wire S3192;
wire S3193;
wire S3194;
wire S3195;
wire S3196;
wire S3197;
wire S3198;
wire S3199;
wire S3200;
wire S3201;
wire S3202;
wire S3203;
wire S3204;
wire S3205;
wire S3206;
wire S3207;
wire S3208;
wire S3209;
wire S3210;
wire S3211;
wire S3212;
wire S3213;
wire S3214;
wire S3215;
wire S3216;
wire S3217;
wire S3218;
wire S3219;
wire S3220;
wire S3221;
wire S3222;
wire S3223;
wire S3224;
wire S3225;
wire S3226;
wire S3227;
wire S3228;
wire S3229;
wire S3230;
wire S3231;
wire S3232;
wire S3233;
wire S3234;
wire S3235;
wire S3236;
wire S3237;
wire S3238;
wire S3239;
wire S3240;
wire S3241;
wire S3242;
wire S3243;
wire S3244;
wire S3245;
wire S3246;
wire S3247;
wire S3248;
wire S3249;
wire S3250;
wire S3251;
wire S3252;
wire S3253;
wire S3254;
wire S3255;
wire S3256;
wire S3257;
wire S3258;
wire S3259;
wire S3260;
wire S3261;
wire S3262;
wire S3263;
wire S3264;
wire S3265;
wire S3266;
wire S3267;
wire S3268;
wire S3269;
wire S3270;
wire S3271;
wire S3272;
wire S3273;
wire S3274;
wire S3275;
wire S3276;
wire S3277;
wire S3278;
wire S3279;
wire S3280;
wire S3281;
wire S3282;
wire S3283;
wire S3284;
wire S3285;
wire S3286;
wire S3287;
wire S3288;
wire S3289;
wire S3290;
wire S3291;
wire S3292;
wire S3293;
wire S3294;
wire S3295;
wire S3296;
wire S3297;
wire S3298;
wire S3299;
wire S3300;
wire S3301;
wire S3302;
wire S3303;
wire S3304;
wire S3305;
wire S3306;
wire S3307;
wire S3308;
wire S3309;
wire S3310;
wire S3311;
wire S3312;
wire S3313;
wire S3314;
wire S3315;
wire S3316;
wire S3317;
wire S3318;
wire S3319;
wire S3320;
wire S3321;
wire S3322;
wire S3323;
wire S3324;
wire S3325;
wire S3326;
wire S3327;
wire S3328;
wire S3329;
wire S3330;
wire S3331;
wire S3332;
wire S3333;
wire S3334;
wire S3335;
wire S3336;
wire S3337;
wire S3338;
wire S3339;
wire S3340;
wire S3341;
wire S3342;
wire S3343;
wire S3344;
wire S3345;
wire S3346;
wire S3347;
wire S3348;
wire S3349;
wire S3350;
wire S3351;
wire S3352;
wire S3353;
wire S3354;
wire S3355;
wire S3356;
wire S3357;
wire S3358;
wire S3359;
wire S3360;
wire S3361;
wire S3362;
wire S3363;
wire S3364;
wire S3365;
wire S3366;
wire S3367;
wire S3368;
wire S3369;
wire S3370;
wire S3371;
wire S3372;
wire S3373;
wire S3374;
wire S3375;
wire S3376;
wire S3377;
wire S3378;
wire S3379;
wire S3380;
wire S3381;
wire S3382;
wire S3383;
wire S3384;
wire S3385;
wire S3386;
wire S3387;
wire S3388;
wire S3389;
wire S3390;
wire S3391;
wire S3392;
wire S3393;
wire S3394;
wire S3395;
wire S3396;
wire S3397;
wire S3398;
wire S3399;
wire S3400;
wire S3401;
wire S3402;
wire S3403;
wire S3404;
wire S3405;
wire S3406;
wire S3407;
wire S3408;
wire S3409;
wire S3410;
wire S3411;
wire S3412;
wire S3413;
wire S3414;
wire S3415;
wire S3416;
wire S3417;
wire S3418;
wire S3419;
wire S3420;
wire S3421;
wire S3422;
wire S3423;
wire S3424;
wire S3425;
wire S3426;
wire S3427;
wire S3428;
wire S3429;
wire S3430;
wire S3431;
wire S3432;
wire S3433;
wire S3434;
wire S3435;
wire S3436;
wire S3437;
wire S3438;
wire S3439;
wire S3440;
wire S3441;
wire S3442;
wire S3443;
wire S3444;
wire S3445;
wire S3446;
wire S3447;
wire S3448;
wire S3449;
wire S3450;
wire S3451;
wire S3452;
wire S3453;
wire S3454;
wire S3455;
wire S3456;
wire S3457;
wire S3458;
wire S3459;
wire S3460;
wire S3461;
wire S3462;
wire S3463;
wire S3464;
wire S3465;
wire S3466;
wire S3467;
wire S3468;
wire S3469;
wire S3470;
wire S3471;
wire S3472;
wire S3473;
wire S3474;
wire S3475;
wire S3476;
wire S3477;
wire S3478;
wire S3479;
wire S3480;
wire S3481;
wire S3482;
wire S3483;
wire S3484;
wire S3485;
wire S3486;
wire S3487;
wire S3488;
wire S3489;
wire S3490;
wire S3491;
wire S3492;
wire S3493;
wire S3494;
wire S3495;
wire S3496;
wire S3497;
wire S3498;
wire S3499;
wire S3500;
wire S3501;
wire S3502;
wire S3503;
wire S3504;
wire S3505;
wire S3506;
wire S3507;
wire S3508;
wire S3509;
wire S3510;
wire S3511;
wire S3512;
wire S3513;
wire S3514;
wire S3515;
wire S3516;
wire S3517;
wire S3518;
wire S3519;
wire S3520;
wire S3521;
wire S3522;
wire S3523;
wire S3524;
wire S3525;
wire S3526;
wire S3527;
wire S3528;
wire S3529;
wire S3530;
wire S3531;
wire S3532;
wire S3533;
wire S3534;
wire S3535;
wire S3536;
wire S3537;
wire S3538;
wire S3539;
wire S3540;
wire S3541;
wire S3542;
wire S3543;
wire S3544;
wire S3545;
wire S3546;
wire S3547;
wire S3548;
wire S3549;
wire S3550;
wire S3551;
wire S3552;
wire S3553;
wire S3554;
wire S3555;
wire S3556;
wire S3557;
wire S3558;
wire S3559;
wire S3560;
wire S3561;
wire S3562;
wire S3563;
wire S3564;
wire S3565;
wire S3566;
wire S3567;
wire S3568;
wire S3569;
wire S3570;
wire S3571;
wire S3572;
wire S3573;
wire S3574;
wire S3575;
wire S3576;
wire S3577;
wire S3578;
wire S3579;
wire S3580;
wire S3581;
wire S3582;
wire S3583;
wire S3584;
wire S3585;
wire S3586;
wire S3587;
wire S3588;
wire S3589;
wire S3590;
wire S3591;
wire S3592;
wire S3593;
wire S3594;
wire S3595;
wire S3596;
wire S3597;
wire S3598;
wire S3599;
wire S3600;
wire S3601;
wire S3602;
wire S3603;
wire S3604;
wire S3605;
wire S3606;
wire S3607;
wire S3608;
wire S3609;
wire S3610;
wire S3611;
wire S3612;
wire S3613;
wire S3614;
wire S3615;
wire S3616;
wire S3617;
wire S3618;
wire S3619;
wire S3620;
wire S3621;
wire S3622;
wire S3623;
wire S3624;
wire S3625;
wire S3626;
wire S3627;
wire S3628;
wire S3629;
wire S3630;
wire S3631;
wire S3632;
wire S3633;
wire S3634;
wire S3635;
wire S3636;
wire S3637;
wire S3638;
wire S3639;
wire S3640;
wire S3641;
wire S3642;
wire S3643;
wire S3644;
wire S3645;
wire S3646;
wire S3647;
wire S3648;
wire S3649;
wire S3650;
wire S3651;
wire S3652;
wire S3653;
wire S3654;
wire S3655;
wire S3656;
wire S3657;
wire S3658;
wire S3659;
wire S3660;
wire S3661;
wire S3662;
wire S3663;
wire S3664;
wire S3665;
wire S3666;
wire S3667;
wire S3668;
wire S3669;
wire S3670;
wire S3671;
wire S3672;
wire S3673;
wire S3674;
wire S3675;
wire S3676;
wire S3677;
wire S3678;
wire S3679;
wire S3680;
wire S3681;
wire S3682;
wire S3683;
wire S3684;
wire S3685;
wire S3686;
wire S3687;
wire S3688;
wire S3689;
wire S3690;
wire S3691;
wire S3692;
wire S3693;
wire S3694;
wire S3695;
wire S3696;
wire S3697;
wire S3698;
wire S3699;
wire S3700;
wire S3701;
wire S3702;
wire S3703;
wire S3704;
wire S3705;
wire S3706;
wire S3707;
wire S3708;
wire S3709;
wire S3710;
wire S3711;
wire S3712;
wire S3713;
wire S3714;
wire S3715;
wire S3716;
wire S3717;
wire S3718;
wire S3719;
wire S3720;
wire S3721;
wire S3722;
wire S3723;
wire S3724;
wire S3725;
wire S3726;
wire S3727;
wire S3728;
wire S3729;
wire S3730;
wire S3731;
wire S3732;
wire S3733;
wire S3734;
wire S3735;
wire S3736;
wire S3737;
wire S3738;
wire S3739;
wire S3740;
wire S3741;
wire S3742;
wire S3743;
wire S3744;
wire S3745;
wire S3746;
wire S3747;
wire S3748;
wire S3749;
wire S3750;
wire S3751;
wire S3752;
wire S3753;
wire S3754;
wire S3755;
wire S3756;
wire S3757;
wire S3758;
wire S3759;
wire S3760;
wire S3761;
wire S3762;
wire S3763;
wire S3764;
wire S3765;
wire S3766;
wire S3767;
wire S3768;
wire S3769;
wire S3770;
wire S3771;
wire S3772;
wire S3773;
wire S3774;
wire S3775;
wire S3776;
wire S3777;
wire S3778;
wire S3779;
wire S3780;
wire S3781;
wire S3782;
wire S3783;
wire S3784;
wire S3785;
wire S3786;
wire S3787;
wire S3788;
wire S3789;
wire S3790;
wire S3791;
wire S3792;
wire S3793;
wire S3794;
wire S3795;
wire S3796;
wire S3797;
wire S3798;
wire S3799;
wire S3800;
wire S3801;
wire S3802;
wire S3803;
wire S3804;
wire S3805;
wire S3806;
wire S3807;
wire S3808;
wire S3809;
wire S3810;
wire S3811;
wire S3812;
wire S3813;
wire S3814;
wire S3815;
wire S3816;
wire S3817;
wire S3818;
wire S3819;
wire S3820;
wire S3821;
wire S3822;
wire S3823;
wire S3824;
wire S3825;
wire S3826;
wire S3827;
wire S3828;
wire S3829;
wire S3830;
wire S3831;
wire S3832;
wire S3833;
wire S3834;
wire S3835;
wire S3836;
wire S3837;
wire S3838;
wire S3839;
wire S3840;
wire S3841;
wire S3842;
wire S3843;
wire S3844;
wire S3845;
wire S3846;
wire S3847;
wire S3848;
wire S3849;
wire S3850;
wire S3851;
wire S3852;
wire S3853;
wire S3854;
wire S3855;
wire S3856;
wire S3857;
wire S3858;
wire S3859;
wire S3860;
wire S3861;
wire S3862;
wire S3863;
wire S3864;
wire S3865;
wire S3866;
wire S3867;
wire S3868;
wire S3869;
wire S3870;
wire S3871;
wire S3872;
wire S3873;
wire S3874;
wire S3875;
wire S3876;
wire S3877;
wire S3878;
wire S3879;
wire S3880;
wire S3881;
wire S3882;
wire S3883;
wire S3884;
wire S3885;
wire S3886;
wire S3887;
wire S3888;
wire S3889;
wire S3890;
wire S3891;
wire S3892;
wire S3893;
wire S3894;
wire S3895;
wire S3896;
wire S3897;
wire S3898;
wire S3899;
wire S3900;
wire S3901;
wire S3902;
wire S3903;
wire S3904;
wire S3905;
wire S3906;
wire S3907;
wire S3908;
wire S3909;
wire S3910;
wire S3911;
wire S3912;
wire S3913;
wire S3914;
wire S3915;
wire S3916;
wire S3917;
wire S3918;
wire S3919;
wire S3920;
wire S3921;
wire S3922;
wire S3923;
wire S3924;
wire S3925;
wire S3926;
wire S3927;
wire S3928;
wire S3929;
wire S3930;
wire S3931;
wire S3932;
wire S3933;
wire S3934;
wire S3935;
wire S3936;
wire S3937;
wire S3938;
wire S3939;
wire S3940;
wire S3941;
wire S3942;
wire S3943;
wire S3944;
wire S3945;
wire S3946;
wire S3947;
wire S3948;
wire S3949;
wire S3950;
wire S3951;
wire S3952;
wire S3953;
wire S3954;
wire S3955;
wire S3956;
wire S3957;
wire S3958;
wire S3959;
wire S3960;
wire S3961;
wire S3962;
wire S3963;
wire S3964;
wire S3965;
wire S3966;
wire S3967;
wire S3968;
wire S3969;
wire S3970;
wire S3971;
wire S3972;
wire S3973;
wire S3974;
wire S3975;
wire S3976;
wire S3977;
wire S3978;
wire S3979;
wire S3980;
wire S3981;
wire S3982;
wire S3983;
wire S3984;
wire S3985;
wire S3986;
wire S3987;
wire S3988;
wire S3989;
wire S3990;
wire S3991;
wire S3992;
wire S3993;
wire S3994;
wire S3995;
wire S3996;
wire S3997;
wire S3998;
wire S3999;
wire S4000;
wire S4001;
wire S4002;
wire S4003;
wire S4004;
wire S4005;
wire S4006;
wire S4007;
wire S4008;
wire S4009;
wire S4010;
wire S4011;
wire S4012;
wire S4013;
wire S4014;
wire S4015;
wire S4016;
wire S4017;
wire S4018;
wire S4019;
wire S4020;
wire S4021;
wire S4022;
wire S4023;
wire S4024;
wire S4025;
wire S4026;
wire S4027;
wire S4028;
wire S4029;
wire S4030;
wire S4031;
wire S4032;
wire S4033;
wire S4034;
wire S4035;
wire S4036;
wire S4037;
wire S4038;
wire S4039;
wire S4040;
wire S4041;
wire S4042;
wire S4043;
wire S4044;
wire S4045;
wire S4046;
wire S4047;
wire S4048;
wire S4049;
wire S4050;
wire S4051;
wire S4052;
wire S4053;
wire S4054;
wire S4055;
wire S4056;
wire S4057;
wire S4058;
wire S4059;
wire S4060;
wire S4061;
wire S4062;
wire S4063;
wire S4064;
wire S4065;
wire S4066;
wire S4067;
wire S4068;
wire S4069;
wire S4070;
wire S4071;
wire S4072;
wire S4073;
wire S4074;
wire S4075;
wire S4076;
wire S4077;
wire S4078;
wire S4079;
wire S4080;
wire S4081;
wire S4082;
wire S4083;
wire S4084;
wire S4085;
wire S4086;
wire S4087;
wire S4088;
wire S4089;
wire S4090;
wire S4091;
wire S4092;
wire S4093;
wire S4094;
wire S4095;
wire S4096;
wire S4097;
wire S4098;
wire S4099;
wire S4100;
wire S4101;
wire S4102;
wire S4103;
wire S4104;
wire S4105;
wire S4106;
wire S4107;
wire S4108;
wire S4109;
wire S4110;
wire S4111;
wire S4112;
wire S4113;
wire S4114;
wire S4115;
wire S4116;
wire S4117;
wire S4118;
wire S4119;
wire S4120;
wire S4121;
wire S4122;
wire S4123;
wire S4124;
wire S4125;
wire S4126;
wire S4127;
wire S4128;
wire S4129;
wire S4130;
wire S4131;
wire S4132;
wire S4133;
wire S4134;
wire S4135;
wire S4136;
wire S4137;
wire S4138;
wire S4139;
wire S4140;
wire S4141;
wire S4142;
wire S4143;
wire S4144;
wire S4145;
wire S4146;
wire S4147;
wire S4148;
wire S4149;
wire S4150;
wire S4151;
wire S4152;
wire S4153;
wire S4154;
wire S4155;
wire S4156;
wire S4157;
wire S4158;
wire S4159;
wire S4160;
wire S4161;
wire S4162;
wire S4163;
wire S4164;
wire S4165;
wire S4166;
wire S4167;
wire S4168;
wire S4169;
wire S4170;
wire S4171;
wire S4172;
wire S4173;
wire S4174;
wire S4175;
wire S4176;
wire S4177;
wire S4178;
wire S4179;
wire S4180;
wire S4181;
wire S4182;
wire S4183;
wire S4184;
wire S4185;
wire S4186;
wire S4187;
wire S4188;
wire S4189;
wire S4190;
wire S4191;
wire S4192;
wire S4193;
wire S4194;
wire S4195;
wire S4196;
wire S4197;
wire S4198;
wire S4199;
wire S4200;
wire S4201;
wire S4202;
wire S4203;
wire S4204;
wire S4205;
wire S4206;
wire S4207;
wire S4208;
wire S4209;
wire S4210;
wire S4211;
wire S4212;
wire S4213;
wire S4214;
wire S4215;
wire S4216;
wire S4217;
wire S4218;
wire S4219;
wire S4220;
wire S4221;
wire S4222;
wire S4223;
wire S4224;
wire S4225;
wire S4226;
wire S4227;
wire S4228;
wire S4229;
wire S4230;
wire S4231;
wire S4232;
wire S4233;
wire S4234;
wire S4235;
wire S4236;
wire S4237;
wire S4238;
wire S4239;
wire S4240;
wire S4241;
wire S4242;
wire S4243;
wire S4244;
wire S4245;
wire S4246;
wire S4247;
wire S4248;
wire S4249;
wire S4250;
wire S4251;
wire S4252;
wire S4253;
wire S4254;
wire S4255;
wire S4256;
wire S4257;
wire S4258;
wire S4259;
wire S4260;
wire S4261;
wire S4262;
wire S4263;
wire S4264;
wire S4265;
wire S4266;
wire S4267;
wire S4268;
wire S4269;
wire S4270;
wire S4271;
wire S4272;
wire S4273;
wire S4274;
wire S4275;
wire S4276;
wire S4277;
wire S4278;
wire S4279;
wire S4280;
wire S4281;
wire S4282;
wire S4283;
wire S4284;
wire S4285;
wire S4286;
wire S4287;
wire S4288;
wire S4289;
wire S4290;
wire S4291;
wire S4292;
wire S4293;
wire S4294;
wire S4295;
wire S4296;
wire S4297;
wire S4298;
wire S4299;
wire S4300;
wire S4301;
wire S4302;
wire S4303;
wire S4304;
wire S4305;
wire S4306;
wire S4307;
wire S4308;
wire S4309;
wire S4310;
wire S4311;
wire S4312;
wire S4313;
wire S4314;
wire S4315;
wire S4316;
wire S4317;
wire S4318;
wire S4319;
wire S4320;
wire S4321;
wire S4322;
wire S4323;
wire S4324;
wire S4325;
wire S4326;
wire S4327;
wire S4328;
wire S4329;
wire S4330;
wire S4331;
wire S4332;
wire S4333;
wire S4334;
wire S4335;
wire S4336;
wire S4337;
wire S4338;
wire S4339;
wire S4340;
wire S4341;
wire S4342;
wire S4343;
wire S4344;
wire S4345;
wire S4346;
wire S4347;
wire S4348;
wire S4349;
wire S4350;
wire S4351;
wire S4352;
wire S4353;
wire S4354;
wire S4355;
wire S4356;
wire S4357;
wire S4358;
wire S4359;
wire S4360;
wire S4361;
wire S4362;
wire S4363;
wire S4364;
wire S4365;
wire S4366;
wire S4367;
wire S4368;
wire S4369;
wire S4370;
wire S4371;
wire S4372;
wire S4373;
wire S4374;
wire S4375;
wire S4376;
wire S4377;
wire S4378;
wire S4379;
wire S4380;
wire S4381;
wire S4382;
wire S4383;
wire S4384;
wire S4385;
wire S4386;
wire S4387;
wire S4388;
wire S4389;
wire S4390;
wire S4391;
wire S4392;
wire S4393;
wire S4394;
wire S4395;
wire S4396;
wire S4397;
wire S4398;
wire S4399;
wire S4400;
wire S4401;
wire S4402;
wire S4403;
wire S4404;
wire S4405;
wire S4406;
wire S4407;
wire S4408;
wire S4409;
wire S4410;
wire S4411;
wire S4412;
wire S4413;
wire S4414;
wire S4415;
wire S4416;
wire S4417;
wire S4418;
wire S4419;
wire S4420;
wire S4421;
wire S4422;
wire S4423;
wire S4424;
wire S4425;
wire S4426;
wire S4427;
wire S4428;
wire S4429;
wire S4430;
wire S4431;
wire S4432;
wire S4433;
wire S4434;
wire S4435;
wire S4436;
wire S4437;
wire S4438;
wire S4439;
wire S4440;
wire S4441;
wire S4442;
wire S4443;
wire S4444;
wire S4445;
wire S4446;
wire S4447;
wire S4448;
wire S4449;
wire S4450;
wire S4451;
wire S4452;
wire S4453;
wire S4454;
wire S4455;
wire S4456;
wire S4457;
wire S4458;
wire S4459;
wire S4460;
wire S4461;
wire S4462;
wire S4463;
wire S4464;
wire S4465;
wire S4466;
wire S4467;
wire S4468;
wire S4469;
wire S4470;
wire S4471;
wire S4472;
wire S4473;
wire S4474;
wire S4475;
wire S4476;
wire S4477;
wire S4478;
wire S4479;
wire S4480;
wire S4481;
wire S4482;
wire S4483;
wire S4484;
wire S4485;
wire S4486;
wire S4487;
wire S4488;
wire S4489;
wire S4490;
wire S4491;
wire S4492;
wire S4493;
wire S4494;
wire S4495;
wire S4496;
wire S4497;
wire S4498;
wire S4499;
wire S4500;
wire S4501;
wire S4502;
wire S4503;
wire S4504;
wire S4505;
wire S4506;
wire S4507;
wire S4508;
wire S4509;
wire S4510;
wire S4511;
wire S4512;
wire S4513;
wire S4514;
wire S4515;
wire S4516;
wire S4517;
wire S4518;
wire S4519;
wire S4520;
wire S4521;
wire S4522;
wire S4523;
wire S4524;
wire S4525;
wire S4526;
wire S4527;
wire S4528;
wire S4529;
wire S4530;
wire S4531;
wire S4532;
wire S4533;
wire S4534;
wire S4535;
wire S4536;
wire S4537;
wire S4538;
wire S4539;
wire S4540;
wire S4541;
wire S4542;
wire S4543;
wire S4544;
wire S4545;
wire S4546;
wire S4547;
wire S4548;
wire S4549;
wire S4550;
wire S4551;
wire S4552;
wire S4553;
wire S4554;
wire S4555;
wire S4556;
wire S4557;
wire S4558;
wire S4559;
wire S4560;
wire S4561;
wire S4562;
wire S4563;
wire S4564;
wire S4565;
wire S4566;
wire S4567;
wire S4568;
wire S4569;
wire S4570;
wire S4571;
wire S4572;
wire S4573;
wire S4574;
wire S4575;
wire S4576;
wire S4577;
wire S4578;
wire S4579;
wire S4580;
wire S4581;
wire S4582;
wire S4583;
wire S4584;
wire S4585;
wire S4586;
wire S4587;
wire S4588;
wire S4589;
wire S4590;
wire S4591;
wire S4592;
wire S4593;
wire S4594;
wire S4595;
wire S4596;
wire S4597;
wire S4598;
wire S4599;
wire S4600;
wire S4601;
wire S4602;
wire S4603;
wire S4604;
wire S4605;
wire S4606;
wire S4607;
wire S4608;
wire S4609;
wire S4610;
wire S4611;
wire S4612;
wire S4613;
wire S4614;
wire S4615;
wire S4616;
wire S4617;
wire S4618;
wire S4619;
wire S4620;
wire S4621;
wire S4622;
wire S4623;
wire S4624;
wire S4625;
wire S4626;
wire S4627;
wire S4628;
wire S4629;
wire S4630;
wire S4631;
wire S4632;
wire S4633;
wire S4634;
wire S4635;
wire S4636;
wire S4637;
wire S4638;
wire S4639;
wire S4640;
wire S4641;
wire S4642;
wire S4643;
wire S4644;
wire S4645;
wire S4646;
wire S4647;
wire S4648;
wire S4649;
wire S4650;
wire S4651;
wire S4652;
wire S4653;
wire S4654;
wire S4655;
wire S4656;
wire S4657;
wire S4658;
wire S4659;
wire S4660;
wire S4661;
wire S4662;
wire S4663;
wire S4664;
wire S4665;
wire S4666;
wire S4667;
wire S4668;
wire S4669;
wire S4670;
wire S4671;
wire S4672;
wire S4673;
wire S4674;
wire S4675;
wire S4676;
wire S4677;
wire S4678;
wire S4679;
wire S4680;
wire S4681;
wire S4682;
wire S4683;
wire S4684;
wire S4685;
wire S4686;
wire S4687;
wire S4688;
wire S4689;
wire S4690;
wire S4691;
wire S4692;
wire S4693;
wire S4694;
wire S4695;
wire S4696;
wire S4697;
wire S4698;
wire S4699;
wire S4700;
wire S4701;
wire S4702;
wire S4703;
wire S4704;
wire S4705;
wire S4706;
wire S4707;
wire S4708;
wire S4709;
wire S4710;
wire S4711;
wire S4712;
wire S4713;
wire S4714;
wire S4715;
wire S4716;
wire S4717;
wire S4718;
wire S4719;
wire S4720;
wire S4721;
wire S4722;
wire S4723;
wire S4724;
wire S4725;
wire S4726;
wire S4727;
wire S4728;
wire S4729;
wire S4730;
wire S4731;
wire S4732;
wire S4733;
wire S4734;
wire S4735;
wire S4736;
wire S4737;
wire S4738;
wire S4739;
wire S4740;
wire S4741;
wire S4742;
wire S4743;
wire S4744;
wire S4745;
wire S4746;
wire S4747;
wire S4748;
wire S4749;
wire S4750;
wire S4751;
wire S4752;
wire S4753;
wire S4754;
wire S4755;
wire S4756;
wire S4757;
wire S4758;
wire S4759;
wire S4760;
wire S4761;
wire S4762;
wire S4763;
wire S4764;
wire S4765;
wire S4766;
wire S4767;
wire S4768;
wire S4769;
wire S4770;
wire S4771;
wire S4772;
wire S4773;
wire S4774;
wire S4775;
wire S4776;
wire S4777;
wire S4778;
wire S4779;
wire S4780;
wire S4781;
wire S4782;
wire S4783;
wire S4784;
wire S4785;
wire S4786;
wire S4787;
wire S4788;
wire S4789;
wire S4790;
wire S4791;
wire S4792;
wire S4793;
wire S4794;
wire S4795;
wire S4796;
wire S4797;
wire S4798;
wire S4799;
wire S4800;
wire S4801;
wire S4802;
wire S4803;
wire S4804;
wire S4805;
wire S4806;
wire S4807;
wire S4808;
wire S4809;
wire S4810;
wire S4811;
wire S4812;
wire S4813;
wire S4814;
wire S4815;
wire S4816;
wire S4817;
wire S4818;
wire S4819;
wire S4820;
wire S4821;
wire S4822;
wire S4823;
wire S4824;
wire S4825;
wire S4826;
wire S4827;
wire S4828;
wire S4829;
wire S4830;
wire S4831;
wire S4832;
wire S4833;
wire S4834;
wire S4835;
wire S4836;
wire S4837;
wire S4838;
wire S4839;
wire S4840;
wire S4841;
wire S4842;
wire S4843;
wire S4844;
wire S4845;
wire S4846;
wire S4847;
wire S4848;
wire S4849;
wire S4850;
wire S4851;
wire S4852;
wire S4853;
wire S4854;
wire S4855;
wire S4856;
wire S4857;
wire S4858;
wire S4859;
wire S4860;
wire S4861;
wire S4862;
wire S4863;
wire S4864;
wire S4865;
wire S4866;
wire S4867;
wire S4868;
wire S4869;
wire S4870;
wire S4871;
wire S4872;
wire S4873;
wire S4874;
wire S4875;
wire S4876;
wire S4877;
wire S4878;
wire S4879;
wire S4880;
wire S4881;
wire S4882;
wire S4883;
wire S4884;
wire S4885;
wire S4886;
wire S4887;
wire S4888;
wire S4889;
wire S4890;
wire S4891;
wire S4892;
wire S4893;
wire S4894;
wire S4895;
wire S4896;
wire S4897;
wire S4898;
wire S4899;
wire S4900;
wire S4901;
wire S4902;
wire S4903;
wire S4904;
wire S4905;
wire S4906;
wire S4907;
wire S4908;
wire S4909;
wire S4910;
wire S4911;
wire S4912;
wire S4913;
wire S4914;
wire S4915;
wire S4916;
wire S4917;
wire S4918;
wire S4919;
wire S4920;
wire S4921;
wire S4922;
wire S4923;
wire S4924;
wire S4925;
wire S4926;
wire S4927;
wire S4928;
wire S4929;
wire S4930;
wire S4931;
wire S4932;
wire S4933;
wire S4934;
wire S4935;
wire S4936;
wire S4937;
wire S4938;
wire S4939;
wire S4940;
wire S4941;
wire S4942;
wire S4943;
wire S4944;
wire S4945;
wire S4946;
wire S4947;
wire S4948;
wire S4949;
wire S4950;
wire S4951;
wire S4952;
wire S4953;
wire S4954;
wire S4955;
wire S4956;
wire S4957;
wire S4958;
wire S4959;
wire S4960;
wire S4961;
wire S4962;
wire S4963;
wire S4964;
wire S4965;
wire S4966;
wire S4967;
wire S4968;
wire S4969;
wire S4970;
wire S4971;
wire S4972;
wire S4973;
wire S4974;
wire S4975;
wire S4976;
wire S4977;
wire S4978;
wire S4979;
wire S4980;
wire S4981;
wire S4982;
wire S4983;
wire S4984;
wire S4985;
wire S4986;
wire S4987;
wire S4988;
wire S4989;
wire S4990;
wire S4991;
wire S4992;
wire S4993;
wire S4994;
wire S4995;
wire S4996;
wire S4997;
wire S4998;
wire S4999;
wire S5000;
wire S5001;
wire S5002;
wire S5003;
wire S5004;
wire S5005;
wire S5006;
wire S5007;
wire S5008;
wire S5009;
wire S5010;
wire S5011;
wire S5012;
wire S5013;
wire S5014;
wire S5015;
wire S5016;
wire S5017;
wire S5018;
wire S5019;
wire S5020;
wire S5021;
wire S5022;
wire S5023;
wire S5024;
wire S5025;
wire S5026;
wire S5027;
wire S5028;
wire S5029;
wire S5030;
wire S5031;
wire S5032;
wire S5033;
wire S5034;
wire S5035;
wire S5036;
wire S5037;
wire S5038;
wire S5039;
wire S5040;
wire S5041;
wire S5042;
wire S5043;
wire S5044;
wire S5045;
wire S5046;
wire S5047;
wire S5048;
wire S5049;
wire S5050;
wire S5051;
wire S5052;
wire S5053;
wire S5054;
wire S5055;
wire S5056;
wire S5057;
wire S5058;
wire S5059;
wire S5060;
wire S5061;
wire S5062;
wire S5063;
wire S5064;
wire S5065;
wire S5066;
wire S5067;
wire S5068;
wire S5069;
wire S5070;
wire S5071;
wire S5072;
wire S5073;
wire S5074;
wire S5075;
wire S5076;
wire S5077;
wire S5078;
wire S5079;
wire S5080;
wire S5081;
wire S5082;
wire S5083;
wire S5084;
wire S5085;
wire S5086;
wire S5087;
wire S5088;
wire S5089;
wire S5090;
wire S5091;
wire S5092;
wire S5093;
wire S5094;
wire S5095;
wire S5096;
wire S5097;
wire S5098;
wire S5099;
wire S5100;
wire S5101;
wire S5102;
wire S5103;
wire S5104;
wire S5105;
wire S5106;
wire S5107;
wire S5108;
wire S5109;
wire S5110;
wire S5111;
wire S5112;
wire S5113;
wire S5114;
wire S5115;
wire S5116;
wire S5117;
wire S5118;
wire S5119;
wire S5120;
wire S5121;
wire S5122;
wire S5123;
wire S5124;
wire S5125;
wire S5126;
wire S5127;
wire S5128;
wire S5129;
wire S5130;
wire S5131;
wire S5132;
wire S5133;
wire S5134;
wire S5135;
wire S5136;
wire S5137;
wire S5138;
wire S5139;
wire S5140;
wire S5141;
wire S5142;
wire S5143;
wire S5144;
wire S5145;
wire S5146;
wire S5147;
wire S5148;
wire S5149;
wire S5150;
wire S5151;
wire S5152;
wire S5153;
wire S5154;
wire S5155;
wire S5156;
wire S5157;
wire S5158;
wire S5159;
wire S5160;
wire S5161;
wire S5162;
wire S5163;
wire S5164;
wire S5165;
wire S5166;
wire S5167;
wire S5168;
wire S5169;
wire S5170;
wire S5171;
wire S5172;
wire S5173;
wire S5174;
wire S5175;
wire S5176;
wire S5177;
wire S5178;
wire S5179;
wire S5180;
wire S5181;
wire S5182;
wire S5183;
wire S5184;
wire S5185;
wire S5186;
wire S5187;
wire S5188;
wire S5189;
wire S5190;
wire S5191;
wire S5192;
wire S5193;
wire S5194;
wire S5195;
wire S5196;
wire S5197;
wire S5198;
wire S5199;
wire S5200;
wire S5201;
wire S5202;
wire S5203;
wire S5204;
wire S5205;
wire S5206;
wire S5207;
wire S5208;
wire S5209;
wire S5210;
wire S5211;
wire S5212;
wire S5213;
wire S5214;
wire S5215;
wire S5216;
wire S5217;
wire S5218;
wire S5219;
wire S5220;
wire S5221;
wire S5222;
wire S5223;
wire S5224;
wire S5225;
wire S5226;
wire S5227;
wire S5228;
wire S5229;
wire S5230;
wire S5231;
wire S5232;
wire S5233;
wire S5234;
wire S5235;
wire S5236;
wire S5237;
wire S5238;
wire S5239;
wire S5240;
wire S5241;
wire S5242;
wire S5243;
wire S5244;
wire S5245;
wire S5246;
wire S5247;
wire S5248;
wire S5249;
wire S5250;
wire S5251;
wire S5252;
wire S5253;
wire S5254;
wire S5255;
wire S5256;
wire S5257;
wire S5258;
wire S5259;
wire S5260;
wire S5261;
wire S5262;
wire S5263;
wire S5264;
wire S5265;
wire S5266;
wire S5267;
wire S5268;
wire S5269;
wire S5270;
wire S5271;
wire S5272;
wire S5273;
wire S5274;
wire S5275;
wire S5276;
wire S5277;
wire S5278;
wire S5279;
wire S5280;
wire S5281;
wire S5282;
wire S5283;
wire S5284;
wire S5285;
wire S5286;
wire S5287;
wire S5288;
wire S5289;
wire S5290;
wire S5291;
wire S5292;
wire S5293;
wire S5294;
wire S5295;
wire S5296;
wire S5297;
wire S5298;
wire S5299;
wire S5300;
wire S5301;
wire S5302;
wire S5303;
wire S5304;
wire S5305;
wire S5306;
wire S5307;
wire S5308;
wire S5309;
wire S5310;
wire S5311;
wire S5312;
wire S5313;
wire S5314;
wire S5315;
wire S5316;
wire S5317;
wire S5318;
wire S5319;
wire S5320;
wire S5321;
wire S5322;
wire S5323;
wire S5324;
wire S5325;
wire S5326;
wire S5327;
wire S5328;
wire S5329;
wire S5330;
wire S5331;
wire S5332;
wire S5333;
wire S5334;
wire S5335;
wire S5336;
wire S5337;
wire S5338;
wire S5339;
wire S5340;
wire S5341;
wire S5342;
wire S5343;
wire S5344;
wire S5345;
wire S5346;
wire S5347;
wire S5348;
wire S5349;
wire S5350;
wire S5351;
wire S5352;
wire S5353;
wire S5354;
wire S5355;
wire S5356;
wire S5357;
wire S5358;
wire S5359;
wire S5360;
wire S5361;
wire S5362;
wire S5363;
wire S5364;
wire S5365;
wire S5366;
wire S5367;
wire S5368;
wire S5369;
wire S5370;
wire S5371;
wire S5372;
wire S5373;
wire S5374;
wire S5375;
wire S5376;
wire S5377;
wire S5378;
wire S5379;
wire S5380;
wire S5381;
wire S5382;
wire S5383;
wire S5384;
wire S5385;
wire S5386;
wire S5387;
wire S5388;
wire S5389;
wire S5390;
wire S5391;
wire S5392;
wire S5393;
wire S5394;
wire S5395;
wire S5396;
wire S5397;
wire S5398;
wire S5399;
wire S5400;
wire S5401;
wire S5402;
wire S5403;
wire S5404;
wire S5405;
wire S5406;
wire S5407;
wire S5408;
wire S5409;
wire S5410;
wire S5411;
wire S5412;
wire S5413;
wire S5414;
wire S5415;
wire S5416;
wire S5417;
wire S5418;
wire S5419;
wire S5420;
wire S5421;
wire S5422;
wire S5423;
wire S5424;
wire S5425;
wire S5426;
wire S5427;
wire S5428;
wire S5429;
wire S5430;
wire S5431;
wire S5432;
wire S5433;
wire S5434;
wire S5435;
wire S5436;
wire S5437;
wire S5438;
wire S5439;
wire S5440;
wire S5441;
wire S5442;
wire S5443;
wire S5444;
wire S5445;
wire S5446;
wire S5447;
wire S5448;
wire S5449;
wire S5450;
wire S5451;
wire S5452;
wire S5453;
wire S5454;
wire S5455;
wire S5456;
wire S5457;
wire S5458;
wire S5459;
wire S5460;
wire S5461;
wire S5462;
wire S5463;
wire S5464;
wire S5465;
wire S5466;
wire S5467;
wire S5468;
wire S5469;
wire S5470;
wire S5471;
wire S5472;
wire S5473;
wire S5474;
wire S5475;
wire S5476;
wire S5477;
wire S5478;
wire S5479;
wire S5480;
wire S5481;
wire S5482;
wire S5483;
wire S5484;
wire S5485;
wire S5486;
wire S5487;
wire S5488;
wire S5489;
wire S5490;
wire S5491;
wire S5492;
wire S5493;
wire S5494;
wire S5495;
wire S5496;
wire S5497;
wire S5498;
wire S5499;
wire S5500;
wire S5501;
wire S5502;
wire S5503;
wire S5504;
wire S5505;
wire S5506;
wire S5507;
wire S5508;
wire S5509;
wire S5510;
wire S5511;
wire S5512;
wire S5513;
wire S5514;
wire S5515;
wire S5516;
wire S5517;
wire S5518;
wire S5519;
wire S5520;
wire S5521;
wire S5522;
wire S5523;
wire S5524;
wire S5525;
wire S5526;
wire S5527;
wire S5528;
wire S5529;
wire S5530;
wire S5531;
wire S5532;
wire S5533;
wire S5534;
wire S5535;
wire S5536;
wire S5537;
wire S5538;
wire S5539;
wire S5540;
wire S5541;
wire S5542;
wire S5543;
wire S5544;
wire S5545;
wire S5546;
wire S5547;
wire S5548;
wire S5549;
wire S5550;
wire S5551;
wire S5552;
wire S5553;
wire S5554;
wire S5555;
wire S5556;
wire S5557;
wire S5558;
wire S5559;
wire S5560;
wire S5561;
wire S5562;
wire S5563;
wire S5564;
wire S5565;
wire S5566;
wire S5567;
wire S5568;
wire S5569;
wire S5570;
wire S5571;
wire S5572;
wire S5573;
wire S5574;
wire S5575;
wire S5576;
wire S5577;
wire S5578;
wire S5579;
wire S5580;
wire S5581;
wire S5582;
wire S5583;
wire S5584;
wire S5585;
wire S5586;
wire S5587;
wire S5588;
wire S5589;
wire S5590;
wire S5591;
wire S5592;
wire S5593;
wire S5594;
wire S5595;
wire S5596;
wire S5597;
wire S5598;
wire S5599;
wire S5600;
wire S5601;
wire S5602;
wire S5603;
wire S5604;
wire S5605;
wire S5606;
wire S5607;
wire S5608;
wire S5609;
wire S5610;
wire S5611;
wire S5612;
wire S5613;
wire S5614;
wire S5615;
wire S5616;
wire S5617;
wire S5618;
wire S5619;
wire S5620;
wire S5621;
wire S5622;
wire S5623;
wire S5624;
wire S5625;
wire S5626;
wire S5627;
wire S5628;
wire S5629;
wire S5630;
wire S5631;
wire S5632;
wire S5633;
wire S5634;
wire S5635;
wire S5636;
wire S5637;
wire S5638;
wire S5639;
wire S5640;
wire S5641;
wire S5642;
wire S5643;
wire S5644;
wire S5645;
wire S5646;
wire S5647;
wire S5648;
wire S5649;
wire S5650;
wire S5651;
wire S5652;
wire S5653;
wire S5654;
wire S5655;
wire S5656;
wire S5657;
wire S5658;
wire S5659;
wire S5660;
wire S5661;
wire S5662;
wire S5663;
wire S5664;
wire S5665;
wire S5666;
wire S5667;
wire S5668;
wire S5669;
wire S5670;
wire S5671;
wire S5672;
wire S5673;
wire S5674;
wire S5675;
wire S5676;
wire S5677;
wire S5678;
wire S5679;
wire S5680;
wire S5681;
wire S5682;
wire S5683;
wire S5684;
wire S5685;
wire S5686;
wire S5687;
wire S5688;
wire S5689;
wire S5690;
wire S5691;
wire S5692;
wire S5693;
wire S5694;
wire S5695;
wire S5696;
wire S5697;
wire S5698;
wire S5699;
wire S5700;
wire S5701;
wire S5702;
wire S5703;
wire S5704;
wire S5705;
wire S5706;
wire S5707;
wire S5708;
wire S5709;
wire S5710;
wire S5711;
wire S5712;
wire S5713;
wire S5714;
wire S5715;
wire S5716;
wire S5717;
wire S5718;
wire S5719;
wire S5720;
wire S5721;
wire S5722;
wire S5723;
wire S5724;
wire S5725;
wire S5726;
wire S5727;
wire S5728;
wire S5729;
wire S5730;
wire S5731;
wire S5732;
wire S5733;
wire S5734;
wire S5735;
wire S5736;
wire S5737;
wire S5738;
wire S5739;
wire S5740;
wire S5741;
wire S5742;
wire S5743;
wire S5744;
wire S5745;
wire S5746;
wire S5747;
wire S5748;
wire S5749;
wire S5750;
wire S5751;
wire S5752;
wire S5753;
wire S5754;
wire S5755;
wire S5756;
wire S5757;
wire S5758;
wire S5759;
wire S5760;
wire S5761;
wire S5762;
wire S5763;
wire S5764;
wire S5765;
wire S5766;
wire S5767;
wire S5768;
wire S5769;
wire S5770;
wire S5771;
wire S5772;
wire S5773;
wire S5774;
wire S5775;
wire S5776;
wire S5777;
wire S5778;
wire S5779;
wire S5780;
wire S5781;
wire S5782;
wire S5783;
wire S5784;
wire S5785;
wire S5786;
wire S5787;
wire S5788;
wire S5789;
wire S5790;
wire S5791;
wire S5792;
wire S5793;
wire S5794;
wire S5795;
wire S5796;
wire S5797;
wire S5798;
wire S5799;
wire S5800;
wire S5801;
wire S5802;
wire S5803;
wire S5804;
wire S5805;
wire S5806;
wire S5807;
wire S5808;
wire S5809;
wire S5810;
wire S5811;
wire S5812;
wire S5813;
wire S5814;
wire S5815;
wire S5816;
wire S5817;
wire S5818;
wire S5819;
wire S5820;
wire S5821;
wire S5822;
wire S5823;
wire S5824;
wire S5825;
wire S5826;
wire S5827;
wire S5828;
wire S5829;
wire S5830;
wire S5831;
wire S5832;
wire S5833;
wire S5834;
wire S5835;
wire S5836;
wire S5837;
wire S5838;
wire S5839;
wire S5840;
wire S5841;
wire S5842;
wire S5843;
wire S5844;
wire S5845;
wire S5846;
wire S5847;
wire S5848;
wire S5849;
wire S5850;
wire S5851;
wire S5852;
wire S5853;
wire S5854;
wire S5855;
wire S5856;
wire S5857;
wire S5858;
wire S5859;
wire S5860;
wire S5861;
wire S5862;
wire S5863;
wire S5864;
wire S5865;
wire S5866;
wire S5867;
wire S5868;
wire S5869;
wire S5870;
wire S5871;
wire S5872;
wire S5873;
wire S5874;
wire S5875;
wire S5876;
wire S5877;
wire S5878;
wire S5879;
wire S5880;
wire S5881;
wire S5882;
wire S5883;
wire S5884;
wire S5885;
wire S5886;
wire S5887;
wire S5888;
wire S5889;
wire S5890;
wire S5891;
wire S5892;
wire S5893;
wire S5894;
wire S5895;
wire S5896;
wire S5897;
wire S5898;
wire S5899;
wire S5900;
wire S5901;
wire S5902;
wire S5903;
wire S5904;
wire S5905;
wire S5906;
wire S5907;
wire S5908;
wire S5909;
wire S5910;
wire S5911;
wire S5912;
wire S5913;
wire S5914;
wire S5915;
wire S5916;
wire S5917;
wire S5918;
wire S5919;
wire S5920;
wire S5921;
wire S5922;
wire S5923;
wire S5924;
wire S5925;
wire S5926;
wire S5927;
wire S5928;
wire S5929;
wire S5930;
wire S5931;
wire S5932;
wire S5933;
wire S5934;
wire S5935;
wire S5936;
wire S5937;
wire S5938;
wire S5939;
wire S5940;
wire S5941;
wire S5942;
wire S5943;
wire S5944;
wire S5945;
wire S5946;
wire S5947;
wire S5948;
wire S5949;
wire S5950;
wire S5951;
wire S5952;
wire S5953;
wire S5954;
wire S5955;
wire S5956;
wire S5957;
wire S5958;
wire S5959;
wire S5960;
wire S5961;
wire S5962;
wire S5963;
wire S5964;
wire S5965;
wire S5966;
wire S5967;
wire S5968;
wire S5969;
wire S5970;
wire S5971;
wire S5972;
wire S5973;
wire S5974;
wire S5975;
wire S5976;
wire S5977;
wire S5978;
wire S5979;
wire S5980;
wire S5981;
wire S5982;
wire S5983;
wire S5984;
wire S5985;
wire S5986;
wire S5987;
wire S5988;
wire S5989;
wire S5990;
wire S5991;
wire S5992;
wire S5993;
wire S5994;
wire S5995;
wire S5996;
wire S5997;
wire S5998;
wire S5999;
wire S6000;
wire S6001;
wire S6002;
wire S6003;
wire S6004;
wire S6005;
wire S6006;
wire S6007;
wire S6008;
wire S6009;
wire S6010;
wire S6011;
wire S6012;
wire S6013;
wire S6014;
wire S6015;
wire S6016;
wire S6017;
wire S6018;
wire S6019;
wire S6020;
wire S6021;
wire S6022;
wire S6023;
wire S6024;
wire S6025;
wire S6026;
wire S6027;
wire S6028;
wire S6029;
wire S6030;
wire S6031;
wire S6032;
wire S6033;
wire S6034;
wire S6035;
wire S6036;
wire S6037;
wire S6038;
wire S6039;
wire S6040;
wire S6041;
wire S6042;
wire S6043;
wire S6044;
wire S6045;
wire S6046;
wire S6047;
wire S6048;
wire S6049;
wire S6050;
wire S6051;
wire S6052;
wire S6053;
wire S6054;
wire S6055;
wire S6056;
wire S6057;
wire S6058;
wire S6059;
wire S6060;
wire S6061;
wire S6062;
wire S6063;
wire S6064;
wire S6065;
wire S6066;
wire S6067;
wire S6068;
wire S6069;
wire S6070;
wire S6071;
wire S6072;
wire S6073;
wire S6074;
wire S6075;
wire S6076;
wire S6077;
wire S6078;
wire S6079;
wire S6080;
wire S6081;
wire S6082;
wire S6083;
wire S6084;
wire S6085;
wire S6086;
wire S6087;
wire S6088;
wire S6089;
wire S6090;
wire S6091;
wire S6092;
wire S6093;
wire S6094;
wire S6095;
wire S6096;
wire S6097;
wire S6098;
wire S6099;
wire S6100;
wire S6101;
wire S6102;
wire S6103;
wire S6104;
wire S6105;
wire S6106;
wire S6107;
wire S6108;
wire S6109;
wire S6110;
wire S6111;
wire S6112;
wire S6113;
wire S6114;
wire S6115;
wire S6116;
wire S6117;
wire S6118;
wire S6119;
wire S6120;
wire S6121;
wire S6122;
wire S6123;
wire S6124;
wire S6125;
wire S6126;
wire S6127;
wire S6128;
wire S6129;
wire S6130;
wire S6131;
wire S6132;
wire S6133;
wire S6134;
wire S6135;
wire S6136;
wire S6137;
wire S6138;
wire S6139;
wire S6140;
wire S6141;
wire S6142;
wire S6143;
wire S6144;
wire S6145;
wire S6146;
wire S6147;
wire S6148;
wire S6149;
wire S6150;
wire S6151;
wire S6152;
wire S6153;
wire S6154;
wire S6155;
wire S6156;
wire S6157;
wire S6158;
wire S6159;
wire S6160;
wire S6161;
wire S6162;
wire S6163;
wire S6164;
wire S6165;
wire S6166;
wire S6167;
wire S6168;
wire S6169;
wire S6170;
wire S6171;
wire S6172;
wire S6173;
wire S6174;
wire S6175;
wire S6176;
wire S6177;
wire S6178;
wire S6179;
wire S6180;
wire S6181;
wire S6182;
wire S6183;
wire S6184;
wire S6185;
wire S6186;
wire S6187;
wire S6188;
wire S6189;
wire S6190;
wire S6191;
wire S6192;
wire S6193;
wire S6194;
wire S6195;
wire S6196;
wire S6197;
wire S6198;
wire S6199;
wire S6200;
wire S6201;
wire S6202;
wire S6203;
wire S6204;
wire S6205;
wire S6206;
wire S6207;
wire S6208;
wire S6209;
wire S6210;
wire S6211;
wire S6212;
wire S6213;
wire S6214;
wire S6215;
wire S6216;
wire S6217;
wire S6218;
wire S6219;
wire S6220;
wire S6221;
wire S6222;
wire S6223;
wire S6224;
wire S6225;
wire S6226;
wire S6227;
wire S6228;
wire S6229;
wire S6230;
wire S6231;
wire S6232;
wire S6233;
wire S6234;
wire S6235;
wire S6236;
wire S6237;
wire S6238;
wire S6239;
wire S6240;
wire S6241;
wire S6242;
wire S6243;
wire S6244;
wire S6245;
wire S6246;
wire S6247;
wire S6248;
wire S6249;
wire S6250;
wire S6251;
wire S6252;
wire S6253;
wire S6254;
wire S6255;
wire S6256;
wire S6257;
wire S6258;
wire S6259;
wire S6260;
wire S6261;
wire S6262;
wire S6263;
wire S6264;
wire S6265;
wire S6266;
wire S6267;
wire S6268;
wire S6269;
wire S6270;
wire S6271;
wire S6272;
wire S6273;
wire S6274;
wire S6275;
wire S6276;
wire S6277;
wire S6278;
wire S6279;
wire S6280;
wire S6281;
wire S6282;
wire S6283;
wire S6284;
wire S6285;
wire S6286;
wire S6287;
wire S6288;
wire S6289;
wire S6290;
wire S6291;
wire S6292;
wire S6293;
wire S6294;
wire S6295;
wire S6296;
wire S6297;
wire S6298;
wire S6299;
wire S6300;
wire S6301;
wire S6302;
wire S6303;
wire S6304;
wire S6305;
wire S6306;
wire new_controller_1133_S_0;
wire new_controller_1133_Y;
wire new_controller_1423_Y_0;
wire new_controller_1423_Y_1;
wire new_controller_234_B_0;
wire new_controller_407_B_0;
wire new_controller_407_B_2;
wire new_controller_clk;
wire new_controller_fib_0;
wire new_controller_fib_1;
wire new_controller_fib_2;
wire new_controller_fib_3;
wire new_controller_fib_4;
wire new_controller_opcode_2;
wire new_controller_opcode_3;
wire new_controller_opcode_4;
wire new_controller_opcode_5;
wire new_controller_opcode_6;
wire new_controller_opcode_7;
wire new_controller_outflag_0;
wire new_controller_outflag_1;
wire new_controller_outflag_2;
wire new_controller_outflag_3;
wire new_controller_outflag_6;
wire new_controller_outflag_7;
wire new_controller_pstate_0;
wire new_controller_pstate_1;
wire new_controller_readymem;
wire new_controller_rst;
wire new_datapath_addrbus_0;
wire new_datapath_addrbus_10;
wire new_datapath_addrbus_11;
wire new_datapath_addrbus_12;
wire new_datapath_addrbus_13;
wire new_datapath_addrbus_14;
wire new_datapath_addrbus_15;
wire new_datapath_addrbus_1;
wire new_datapath_addrbus_2;
wire new_datapath_addrbus_3;
wire new_datapath_addrbus_4;
wire new_datapath_addrbus_5;
wire new_datapath_addrbus_6;
wire new_datapath_addrbus_7;
wire new_datapath_addrbus_8;
wire new_datapath_addrbus_9;
wire new_datapath_addsubunit_in1_0;
wire new_datapath_addsubunit_in1_10;
wire new_datapath_addsubunit_in1_11;
wire new_datapath_addsubunit_in1_12;
wire new_datapath_addsubunit_in1_13;
wire new_datapath_addsubunit_in1_14;
wire new_datapath_addsubunit_in1_15;
wire new_datapath_addsubunit_in1_1;
wire new_datapath_addsubunit_in1_2;
wire new_datapath_addsubunit_in1_3;
wire new_datapath_addsubunit_in1_4;
wire new_datapath_addsubunit_in1_5;
wire new_datapath_addsubunit_in1_6;
wire new_datapath_addsubunit_in1_7;
wire new_datapath_addsubunit_in1_8;
wire new_datapath_addsubunit_in1_9;
wire new_datapath_adr_outreg_0;
wire new_datapath_adr_outreg_10;
wire new_datapath_adr_outreg_11;
wire new_datapath_adr_outreg_12;
wire new_datapath_adr_outreg_13;
wire new_datapath_adr_outreg_14;
wire new_datapath_adr_outreg_15;
wire new_datapath_adr_outreg_1;
wire new_datapath_adr_outreg_2;
wire new_datapath_adr_outreg_3;
wire new_datapath_adr_outreg_4;
wire new_datapath_adr_outreg_5;
wire new_datapath_adr_outreg_6;
wire new_datapath_adr_outreg_7;
wire new_datapath_adr_outreg_8;
wire new_datapath_adr_outreg_9;
wire new_datapath_databusin_0;
wire new_datapath_databusin_10;
wire new_datapath_databusin_11;
wire new_datapath_databusin_12;
wire new_datapath_databusin_13;
wire new_datapath_databusin_14;
wire new_datapath_databusin_15;
wire new_datapath_databusin_1;
wire new_datapath_databusin_2;
wire new_datapath_databusin_3;
wire new_datapath_databusin_4;
wire new_datapath_databusin_5;
wire new_datapath_databusin_6;
wire new_datapath_databusin_7;
wire new_datapath_databusin_8;
wire new_datapath_databusin_9;
wire new_datapath_indatatrf_0;
wire new_datapath_indatatrf_10;
wire new_datapath_indatatrf_11;
wire new_datapath_indatatrf_12;
wire new_datapath_indatatrf_13;
wire new_datapath_indatatrf_14;
wire new_datapath_indatatrf_15;
wire new_datapath_indatatrf_1;
wire new_datapath_indatatrf_2;
wire new_datapath_indatatrf_3;
wire new_datapath_indatatrf_4;
wire new_datapath_indatatrf_5;
wire new_datapath_indatatrf_6;
wire new_datapath_indatatrf_7;
wire new_datapath_indatatrf_8;
wire new_datapath_indatatrf_9;
wire new_datapath_instruction_0;
wire new_datapath_instruction_1;
wire new_datapath_instruction_2;
wire new_datapath_instruction_3;
wire new_datapath_multdivunit_1697_B_10;
wire new_datapath_multdivunit_1697_B_11;
wire new_datapath_multdivunit_1697_B_12;
wire new_datapath_multdivunit_1697_B_13;
wire new_datapath_multdivunit_1697_B_14;
wire new_datapath_multdivunit_1697_B_15;
wire new_datapath_multdivunit_1697_B_8;
wire new_datapath_multdivunit_1697_B_9;
wire new_datapath_multdivunit_outmdu1_0;
wire new_datapath_multdivunit_outmdu1_10;
wire new_datapath_multdivunit_outmdu1_11;
wire new_datapath_multdivunit_outmdu1_12;
wire new_datapath_multdivunit_outmdu1_13;
wire new_datapath_multdivunit_outmdu1_14;
wire new_datapath_multdivunit_outmdu1_15;
wire new_datapath_multdivunit_outmdu1_1;
wire new_datapath_multdivunit_outmdu1_2;
wire new_datapath_multdivunit_outmdu1_3;
wire new_datapath_multdivunit_outmdu1_4;
wire new_datapath_multdivunit_outmdu1_5;
wire new_datapath_multdivunit_outmdu1_6;
wire new_datapath_multdivunit_outmdu1_7;
wire new_datapath_multdivunit_outmdu1_8;
wire new_datapath_multdivunit_outmdu1_9;
wire new_datapath_multdivunit_outmdu2_0;
wire new_datapath_multdivunit_outmdu2_10;
wire new_datapath_multdivunit_outmdu2_11;
wire new_datapath_multdivunit_outmdu2_12;
wire new_datapath_multdivunit_outmdu2_13;
wire new_datapath_multdivunit_outmdu2_14;
wire new_datapath_multdivunit_outmdu2_15;
wire new_datapath_multdivunit_outmdu2_1;
wire new_datapath_multdivunit_outmdu2_2;
wire new_datapath_multdivunit_outmdu2_3;
wire new_datapath_multdivunit_outmdu2_4;
wire new_datapath_multdivunit_outmdu2_5;
wire new_datapath_multdivunit_outmdu2_6;
wire new_datapath_multdivunit_outmdu2_7;
wire new_datapath_multdivunit_outmdu2_8;
wire new_datapath_multdivunit_outmdu2_9;
wire new_datapath_muxmem_in2_0;
wire new_datapath_muxmem_in2_10;
wire new_datapath_muxmem_in2_11;
wire new_datapath_muxmem_in2_12;
wire new_datapath_muxmem_in2_13;
wire new_datapath_muxmem_in2_14;
wire new_datapath_muxmem_in2_15;
wire new_datapath_muxmem_in2_1;
wire new_datapath_muxmem_in2_2;
wire new_datapath_muxmem_in2_3;
wire new_datapath_muxmem_in2_4;
wire new_datapath_muxmem_in2_5;
wire new_datapath_muxmem_in2_6;
wire new_datapath_muxmem_in2_7;
wire new_datapath_muxmem_in2_8;
wire new_datapath_muxmem_in2_9;
wire new_datapath_muxrd_outmux_0;
wire new_datapath_muxrd_outmux_1;
wire new_datapath_muxrd_outmux_2;
wire new_datapath_muxrd_outmux_3;
wire new_datapath_muxrs1_outmux_0;
wire new_datapath_muxrs1_outmux_1;
wire new_datapath_muxrs1_outmux_2;
wire new_datapath_muxrs1_outmux_3;
wire new_datapath_muxrs2_outmux_0;
wire new_datapath_muxrs2_outmux_1;
wire new_datapath_muxrs2_outmux_2;
wire new_datapath_muxrs2_outmux_3;
wire new_datapath_p1trf_0;
wire new_datapath_p1trf_1;
wire new_datapath_p1trf_2;
wire new_datapath_p1trf_3;
wire new_datapath_p1trf_4;
wire new_datapath_p1trf_5;
wire new_datapath_p1trf_6;
wire new_datapath_p1trf_7;
wire new_datapath_p2trf_0;
wire new_datapath_p2trf_1;
wire new_datapath_p2trf_2;
wire new_datapath_p2trf_3;
wire new_datapath_p2trf_4;
wire new_datapath_p2trf_5;
wire new_datapath_p2trf_6;
wire new_datapath_p2trf_7;
wire new_datapath_shiftunit_1961_A;
wire new_datapath_shiftunit_1979_A;
wire new_datapath_shiftunit_1997_A;
wire new_datapath_shiftunit_2015_A;
wire new_datapath_shiftunit_2033_A;
wire new_datapath_shiftunit_2051_A;
wire new_datapath_shiftunit_2069_A;
wire new_datapath_shiftunit_2087_A;
wire new_datapath_shiftunit_2105_A;
wire new_datapath_shiftunit_2123_A;
wire new_datapath_shiftunit_2141_A;
wire new_datapath_shiftunit_2159_A;
wire new_datapath_shiftunit_2177_A;
wire new_datapath_shiftunit_2195_A;
wire new_datapath_shiftunit_2213_A;
wire new_datapath_shiftunit_2231_A;
wire new_datapath_shiftunit_2265_A;
wire new_datapath_shiftunit_2283_A;
wire new_datapath_shiftunit_2301_A;
wire new_datapath_shiftunit_2319_A;
wire new_datapath_shiftunit_2337_A;
wire new_datapath_shiftunit_2355_A;
wire new_datapath_shiftunit_2373_A;
wire new_datapath_shiftunit_2391_A;
wire new_datapath_shiftunit_2409_A;
wire new_datapath_shiftunit_2427_A;
wire new_datapath_shiftunit_2445_A;
wire new_datapath_shiftunit_2463_A;
wire new_datapath_shiftunit_2481_A;
wire new_datapath_shiftunit_2499_A;
wire new_datapath_shiftunit_2517_A;
wire new_datapath_shiftunit_2534_A;
input clk;
input rst;
input readyMEM;
input [15:0] dataBusIn;input [15:0] p1TRF;input [15:0] p2TRF;output readMM;
output writeMM;
output [15:0] dataBusOut;output [15:0] addrBus;output [3:0] outMuxrs1;output [3:0] outMuxrs2;output [3:0] outMuxrd;output [15:0] inDataTRF;output writeTRF;
output readInst;

notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_0_ (
  .in1({ new_datapath_multdivunit_outmdu2_15 }),
  .out1({ S2581 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1_ (
  .in1({ new_controller_opcode_7 }),
  .out1({ S2592 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2_ (
  .in1({ new_datapath_databusin_15 }),
  .out1({ S2603 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3_ (
  .in1({ new_controller_outflag_7 }),
  .out1({ S2614 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4_ (
  .in1({ new_datapath_muxmem_in2_0 }),
  .out1({ S2625 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5_ (
  .in1({ new_datapath_muxmem_in2_1 }),
  .out1({ S2636 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6_ (
  .in1({ new_datapath_muxmem_in2_2 }),
  .out1({ S2647 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_7_ (
  .in1({ new_datapath_muxmem_in2_3 }),
  .out1({ S2658 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_8_ (
  .in1({ new_datapath_muxmem_in2_4 }),
  .out1({ S2669 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_9_ (
  .in1({ new_datapath_muxmem_in2_5 }),
  .out1({ S2680 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_10_ (
  .in1({ new_datapath_muxmem_in2_6 }),
  .out1({ S2690 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_11_ (
  .in1({ new_datapath_muxmem_in2_7 }),
  .out1({ S2701 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_12_ (
  .in1({ new_datapath_muxmem_in2_8 }),
  .out1({ S2712 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_13_ (
  .in1({ new_datapath_muxmem_in2_9 }),
  .out1({ S2723 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_14_ (
  .in1({ new_datapath_muxmem_in2_10 }),
  .out1({ S2734 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_15_ (
  .in1({ new_datapath_muxmem_in2_11 }),
  .out1({ S2745 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_16_ (
  .in1({ new_datapath_muxmem_in2_12 }),
  .out1({ S2756 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_17_ (
  .in1({ new_datapath_muxmem_in2_13 }),
  .out1({ S2767 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_18_ (
  .in1({ new_datapath_muxmem_in2_14 }),
  .out1({ S2778 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_19_ (
  .in1({ new_datapath_multdivunit_outmdu1_6 }),
  .out1({ S2789 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_20_ (
  .in1({ new_datapath_multdivunit_outmdu2_0 }),
  .out1({ S2800 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_21_ (
  .in1({ new_datapath_multdivunit_outmdu2_1 }),
  .out1({ S2811 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_22_ (
  .in1({ new_datapath_multdivunit_outmdu2_2 }),
  .out1({ S2822 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_23_ (
  .in1({ new_datapath_multdivunit_outmdu2_3 }),
  .out1({ S2832 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_24_ (
  .in1({ new_datapath_multdivunit_outmdu2_4 }),
  .out1({ S2843 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_25_ (
  .in1({ new_datapath_multdivunit_outmdu2_5 }),
  .out1({ S2854 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_26_ (
  .in1({ new_datapath_multdivunit_outmdu2_6 }),
  .out1({ S2865 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_27_ (
  .in1({ new_datapath_multdivunit_outmdu2_7 }),
  .out1({ S2876 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_28_ (
  .in1({ new_datapath_multdivunit_outmdu2_8 }),
  .out1({ S2887 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_29_ (
  .in1({ new_datapath_multdivunit_outmdu2_9 }),
  .out1({ S2898 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_30_ (
  .in1({ new_datapath_multdivunit_outmdu2_10 }),
  .out1({ S2909 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_31_ (
  .in1({ new_datapath_multdivunit_outmdu2_11 }),
  .out1({ S2920 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_32_ (
  .in1({ new_datapath_multdivunit_outmdu2_12 }),
  .out1({ S2931 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_33_ (
  .in1({ new_datapath_multdivunit_outmdu2_13 }),
  .out1({ S2942 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_34_ (
  .in1({ new_datapath_multdivunit_outmdu2_14 }),
  .out1({ S2953 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_35_ (
  .in1({ new_datapath_instruction_0 }),
  .out1({ S2964 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_36_ (
  .in1({ new_datapath_instruction_3 }),
  .out1({ S2975 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_37_ (
  .in1({ new_controller_fib_0 }),
  .out1({ S2985 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_38_ (
  .in1({ new_controller_fib_1 }),
  .out1({ S2996 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_39_ (
  .in1({ new_controller_fib_2 }),
  .out1({ S3007 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_40_ (
  .in1({ new_controller_fib_3 }),
  .out1({ S3018 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_41_ (
  .in1({ new_controller_fib_4 }),
  .out1({ S3029 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_42_ (
  .in1({ new_controller_234_B_0 }),
  .out1({ S3040 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_43_ (
  .in1({ new_controller_opcode_2 }),
  .out1({ S3051 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_44_ (
  .in1({ new_controller_opcode_3 }),
  .out1({ S3062 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_45_ (
  .in1({ new_controller_opcode_4 }),
  .out1({ S3073 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_46_ (
  .in1({ new_controller_opcode_5 }),
  .out1({ S3084 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_47_ (
  .in1({ new_controller_opcode_6 }),
  .out1({ S3095 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_48_ (
  .in1({ new_datapath_databusin_14 }),
  .out1({ S3106 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_49_ (
  .in1({ new_controller_407_B_0 }),
  .out1({ S3117 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_50_ (
  .in1({ new_controller_pstate_1 }),
  .out1({ S3128 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_51_ (
  .in1({ new_controller_pstate_0 }),
  .out1({ S3139 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_52_ (
  .in1({ new_datapath_p1trf_0 }),
  .out1({ S3150 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_53_ (
  .in1({ new_datapath_p1trf_1 }),
  .out1({ S3160 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_54_ (
  .in1({ new_datapath_p1trf_2 }),
  .out1({ S3171 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_55_ (
  .in1({ new_datapath_p1trf_3 }),
  .out1({ S3182 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_56_ (
  .in1({ new_datapath_p1trf_4 }),
  .out1({ S3193 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_57_ (
  .in1({ new_datapath_p1trf_5 }),
  .out1({ S3204 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_58_ (
  .in1({ new_datapath_p1trf_6 }),
  .out1({ S3215 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_59_ (
  .in1({ new_datapath_p1trf_7 }),
  .out1({ S3226 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_60_ (
  .in1({ new_datapath_p2trf_0 }),
  .out1({ S3237 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_61_ (
  .in1({ new_datapath_p2trf_1 }),
  .out1({ S3248 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_62_ (
  .in1({ new_datapath_p2trf_2 }),
  .out1({ S3259 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_63_ (
  .in1({ new_datapath_p2trf_3 }),
  .out1({ S3270 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_64_ (
  .in1({ new_datapath_p2trf_4 }),
  .out1({ S3281 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_65_ (
  .in1({ new_datapath_p2trf_5 }),
  .out1({ S3292 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_66_ (
  .in1({ new_datapath_p2trf_6 }),
  .out1({ S3303 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_67_ (
  .in1({ new_datapath_p2trf_7 }),
  .out1({ S3314 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_68_ (
  .in1({ new_datapath_addsubunit_in1_8 }),
  .out1({ S3325 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_69_ (
  .in1({ new_datapath_addsubunit_in1_9 }),
  .out1({ S3336 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_70_ (
  .in1({ new_datapath_addsubunit_in1_10 }),
  .out1({ S3346 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_71_ (
  .in1({ new_datapath_addsubunit_in1_11 }),
  .out1({ S3357 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_72_ (
  .in1({ new_datapath_addsubunit_in1_12 }),
  .out1({ S3368 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_73_ (
  .in1({ new_datapath_addsubunit_in1_13 }),
  .out1({ S3379 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_74_ (
  .in1({ new_datapath_addsubunit_in1_14 }),
  .out1({ S3390 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_75_ (
  .in1({ new_datapath_addsubunit_in1_15 }),
  .out1({ S3401 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_76_ (
  .in1({ new_datapath_multdivunit_1697_B_14 }),
  .out1({ S3412 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_77_ (
  .in1({ new_datapath_multdivunit_1697_B_13 }),
  .out1({ S3423 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_78_ (
  .in1({ new_datapath_multdivunit_1697_B_12 }),
  .out1({ S3434 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_79_ (
  .in1({ new_datapath_multdivunit_1697_B_11 }),
  .out1({ S3445 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_80_ (
  .in1({ new_datapath_multdivunit_1697_B_10 }),
  .out1({ S3456 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_81_ (
  .in1({ new_datapath_multdivunit_1697_B_9 }),
  .out1({ S3467 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_82_ (
  .in1({ new_datapath_multdivunit_1697_B_8 }),
  .out1({ S3478 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_83_ (
  .in1({ new_datapath_shiftunit_1997_A }),
  .out1({ S3489 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_84_ (
  .in1({ new_datapath_shiftunit_2015_A }),
  .out1({ S3500 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_85_ (
  .in1({ new_datapath_shiftunit_2069_A }),
  .out1({ S3511 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_86_ (
  .in1({ new_datapath_shiftunit_2087_A }),
  .out1({ S3522 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_87_ (
  .in1({ new_datapath_shiftunit_2105_A }),
  .out1({ S3533 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_88_ (
  .in1({ new_datapath_shiftunit_2123_A }),
  .out1({ S3544 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_89_ (
  .in1({ new_datapath_shiftunit_2141_A }),
  .out1({ S3554 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_90_ (
  .in1({ new_datapath_shiftunit_2159_A }),
  .out1({ S3565 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_91_ (
  .in1({ new_datapath_shiftunit_2177_A }),
  .out1({ S3576 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_92_ (
  .in1({ new_controller_opcode_6, new_controller_opcode_7 }),
  .out1({ S3587 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_93_ (
  .in1({ S3587 }),
  .out1({ S3598 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_94_ (
  .in1({ S3084, new_controller_opcode_4 }),
  .out1({ S3609 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_95_ (
  .in1({ new_controller_opcode_5, S3073 }),
  .out1({ S3620 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_96_ (
  .in1({ S3598, new_controller_opcode_4 }),
  .out1({ S3631 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_97_ (
  .in1({ S3620, S3598 }),
  .out1({ S3642 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_98_ (
  .in1({ S3609, S3587 }),
  .out1({ S3653 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_99_ (
  .in1({ new_controller_pstate_0, S3128 }),
  .out1({ S3664 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_100_ (
  .in1({ S3664 }),
  .out1({ S3675 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_101_ (
  .in1({ S3653, new_controller_opcode_3 }),
  .out1({ S3686 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_102_ (
  .in1({ S3686 }),
  .out1({ S3697 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_103_ (
  .in1({ S3697, S3675 }),
  .out1({ S3708 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_104_ (
  .in1({ S3686, S3664 }),
  .out1({ S3719 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_105_ (
  .in1({ S3719, new_controller_opcode_2 }),
  .out1({ S6215 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_106_ (
  .in1({ S6215 }),
  .out1({ S3740 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_107_ (
  .in1({ S3719, S3051 }),
  .out1({ S6216 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_108_ (
  .in1({ S3139, new_controller_pstate_1 }),
  .out1({ S3761 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_109_ (
  .in1({ new_controller_pstate_0, S3128 }),
  .out1({ S3771 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_110_ (
  .in1({ new_controller_opcode_6, new_controller_opcode_7 }),
  .out1({ S3782 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_111_ (
  .in1({ S3782 }),
  .out1({ S3793 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_112_ (
  .in1({ S3793, S3631 }),
  .out1({ S3804 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_113_ (
  .in1({ S3084, S3073 }),
  .out1({ S3815 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_114_ (
  .in1({ new_controller_opcode_5, new_controller_opcode_4 }),
  .out1({ S3826 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_115_ (
  .in1({ S3826, S3782 }),
  .out1({ S3837 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_116_ (
  .in1({ S3062, new_controller_opcode_2 }),
  .out1({ S3848 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_117_ (
  .in1({ new_controller_opcode_3, S3051 }),
  .out1({ S3859 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_118_ (
  .in1({ S3837, new_controller_opcode_3 }),
  .out1({ S3870 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_119_ (
  .in1({ S3870, new_controller_opcode_2 }),
  .out1({ S3881 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_120_ (
  .in1({ S3881 }),
  .out1({ S3892 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_121_ (
  .in1({ new_controller_opcode_5, new_controller_opcode_4 }),
  .out1({ S3903 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_122_ (
  .in1({ S3084, S3073 }),
  .out1({ S3914 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_123_ (
  .in1({ S3903, S3804 }),
  .out1({ S3925 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_124_ (
  .in1({ S3925, S3892 }),
  .out1({ S3936 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_125_ (
  .in1({ S3642, new_controller_opcode_3 }),
  .out1({ S3947 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_126_ (
  .in1({ S3859, S3837 }),
  .out1({ S3958 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_127_ (
  .in1({ new_controller_opcode_3, S3051 }),
  .out1({ S3969 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_128_ (
  .in1({ S3969, new_controller_fib_2 }),
  .out1({ S3980 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_129_ (
  .in1({ S3980, S2996 }),
  .out1({ S3990 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_130_ (
  .in1({ S3990, S3958 }),
  .out1({ S4001 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_131_ (
  .in1({ S4001 }),
  .out1({ S4012 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_132_ (
  .in1({ S4012, S3947 }),
  .out1({ S4023 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_133_ (
  .in1({ S4023, S3936 }),
  .out1({ S4034 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_134_ (
  .in1({ S4034, S3771 }),
  .out1({ S4045 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_135_ (
  .in1({ new_controller_opcode_5, S3073 }),
  .out1({ S4056 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_136_ (
  .in1({ S3084, new_controller_opcode_4 }),
  .out1({ S4067 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_137_ (
  .in1({ S4056, S3609 }),
  .out1({ S4078 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_138_ (
  .in1({ S4067, S3620 }),
  .out1({ S4089 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_139_ (
  .in1({ S4078, S3782 }),
  .out1({ S4100 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_140_ (
  .in1({ S4100 }),
  .out1({ S4111 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_141_ (
  .in1({ S4111, S3128 }),
  .out1({ S4122 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_142_ (
  .in1({ S4100, new_controller_pstate_1 }),
  .out1({ S4133 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_143_ (
  .in1({ S4133, S3139 }),
  .out1({ S4144 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_144_ (
  .in1({ S4122, new_controller_pstate_0 }),
  .out1({ S4155 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_145_ (
  .in1({ new_controller_readymem, new_controller_234_B_0 }),
  .out1({ S4166 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_146_ (
  .in1({ S4166 }),
  .out1({ S4177 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_147_ (
  .in1({ S4177, S3708 }),
  .out1({ S4188 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_148_ (
  .in1({ S4188, S4155 }),
  .out1({ S4199 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_149_ (
  .in1({ S4199, S4045 }),
  .out1({ S4210 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_150_ (
  .in1({ S4210, new_datapath_muxmem_in2_15 }),
  .out1({ S4221 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_151_ (
  .in1({ S3761, S3609 }),
  .out1({ S4232 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_152_ (
  .in1({ S4232 }),
  .out1({ S4237 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_153_ (
  .in1({ S3771, S3653 }),
  .out1({ S4238 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_154_ (
  .in1({ S3761, S3642 }),
  .out1({ S4246 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_155_ (
  .in1({ S4246, S3062 }),
  .out1({ S4254 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_156_ (
  .in1({ S4238, new_controller_opcode_3 }),
  .out1({ S4261 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_157_ (
  .in1({ new_controller_opcode_3, new_controller_opcode_2 }),
  .out1({ S4269 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_158_ (
  .in1({ S4269 }),
  .out1({ S4278 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_159_ (
  .in1({ S4269, S4246 }),
  .out1({ S4289 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_160_ (
  .in1({ S4289, new_controller_234_B_0 }),
  .out1({ S4300 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_161_ (
  .in1({ S4269, S4238 }),
  .out1({ S4311 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_162_ (
  .in1({ new_controller_407_B_2, new_controller_fib_0 }),
  .out1({ S4322 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_163_ (
  .in1({ S4322 }),
  .out1({ S4333 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_164_ (
  .in1({ new_controller_407_B_2, new_controller_407_B_0 }),
  .out1({ S4344 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_165_ (
  .in1({ new_controller_fib_2, S2996 }),
  .out1({ S4355 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_166_ (
  .in1({ S4355, S4333 }),
  .out1({ S4366 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_167_ (
  .in1({ S4366, S4344 }),
  .out1({ S4377 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_168_ (
  .in1({ new_controller_fib_1, new_controller_fib_0 }),
  .out1({ S4388 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_169_ (
  .in1({ S4388, new_controller_fib_2 }),
  .out1({ S4399 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_170_ (
  .in1({ S4399 }),
  .out1({ S4410 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_171_ (
  .in1({ new_controller_fib_2, S2985 }),
  .out1({ S4421 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_172_ (
  .in1({ S3007, new_controller_fib_0 }),
  .out1({ S4432 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_173_ (
  .in1({ S4432, new_controller_fib_1 }),
  .out1({ S4443 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_174_ (
  .in1({ S4443, S4410 }),
  .out1({ S4454 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_175_ (
  .in1({ S4454, new_controller_407_B_2 }),
  .out1({ S4465 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_176_ (
  .in1({ S4465, new_controller_407_B_0 }),
  .out1({ S4476 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_177_ (
  .in1({ S4388, S3007 }),
  .out1({ S4487 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_178_ (
  .in1({ S4388, S3117 }),
  .out1({ S4498 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_179_ (
  .in1({ S4498, S4476 }),
  .out1({ S4509 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_180_ (
  .in1({ S4509, S4377 }),
  .out1({ S4519 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_181_ (
  .in1({ S4519 }),
  .out1({ S4530 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_182_ (
  .in1({ S3969, new_controller_234_B_0 }),
  .out1({ S4541 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_183_ (
  .in1({ S3782, S3771 }),
  .out1({ S4552 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_184_ (
  .in1({ S3793, S3761 }),
  .out1({ S4563 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_185_ (
  .in1({ S4563, S3826 }),
  .out1({ S4570 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_186_ (
  .in1({ S3837, S3761 }),
  .out1({ S4578 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_187_ (
  .in1({ S4578, S4541 }),
  .out1({ S4586 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_188_ (
  .in1({ S4586, S4530 }),
  .out1({ S4593 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_189_ (
  .in1({ S4593, S4311 }),
  .out1({ S4602 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_190_ (
  .in1({ S4602, new_datapath_addsubunit_in1_14 }),
  .out1({ S4613 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_191_ (
  .in1({ S4613, S4300 }),
  .out1({ S4621 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_192_ (
  .in1({ S4621, new_datapath_muxmem_in2_14 }),
  .out1({ S4632 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_193_ (
  .in1({ S4632 }),
  .out1({ S4643 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_194_ (
  .in1({ S4621, new_datapath_muxmem_in2_14 }),
  .out1({ S4654 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_195_ (
  .in1({ S4654, S4643 }),
  .out1({ S4665 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_196_ (
  .in1({ S4602, new_datapath_addsubunit_in1_13 }),
  .out1({ S4676 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_197_ (
  .in1({ S4676, S4300 }),
  .out1({ S4686 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_198_ (
  .in1({ S4686, new_datapath_muxmem_in2_13 }),
  .out1({ S4697 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_199_ (
  .in1({ S4697 }),
  .out1({ S4708 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_200_ (
  .in1({ S4686, new_datapath_muxmem_in2_13 }),
  .out1({ S4718 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_201_ (
  .in1({ S4602, new_datapath_addsubunit_in1_12 }),
  .out1({ S4729 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_202_ (
  .in1({ S4729, S4300 }),
  .out1({ S4740 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_203_ (
  .in1({ S4740, new_datapath_muxmem_in2_12 }),
  .out1({ S4750 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_204_ (
  .in1({ S4750 }),
  .out1({ S4761 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_205_ (
  .in1({ S4740, new_datapath_muxmem_in2_12 }),
  .out1({ S4772 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_206_ (
  .in1({ S4772, S4761 }),
  .out1({ S4783 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_207_ (
  .in1({ S4602, new_datapath_addsubunit_in1_11 }),
  .out1({ S4793 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_208_ (
  .in1({ S4793, S4300 }),
  .out1({ S4804 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_209_ (
  .in1({ S4804 }),
  .out1({ S4815 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_210_ (
  .in1({ S4804, new_datapath_muxmem_in2_11 }),
  .out1({ S4825 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_211_ (
  .in1({ S4815, S2745 }),
  .out1({ S4836 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_212_ (
  .in1({ S4602, new_datapath_addsubunit_in1_10 }),
  .out1({ S4847 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_213_ (
  .in1({ S4847, S4300 }),
  .out1({ S4857 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_214_ (
  .in1({ S4857, new_datapath_muxmem_in2_10 }),
  .out1({ S4868 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_215_ (
  .in1({ S4868 }),
  .out1({ S4879 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_216_ (
  .in1({ S4857, new_datapath_muxmem_in2_10 }),
  .out1({ S4890 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_217_ (
  .in1({ S4890, S4879 }),
  .out1({ S4900 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_218_ (
  .in1({ S4602, new_datapath_addsubunit_in1_9 }),
  .out1({ S4911 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_219_ (
  .in1({ S4911, S4300 }),
  .out1({ S4922 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_220_ (
  .in1({ S4922, new_datapath_muxmem_in2_9 }),
  .out1({ S4932 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_221_ (
  .in1({ S4932 }),
  .out1({ S4943 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_222_ (
  .in1({ S4922, new_datapath_muxmem_in2_9 }),
  .out1({ S4954 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_223_ (
  .in1({ S4602, new_datapath_addsubunit_in1_8 }),
  .out1({ S4964 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_224_ (
  .in1({ S4964, S4300 }),
  .out1({ S4975 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_225_ (
  .in1({ S4975, new_datapath_muxmem_in2_8 }),
  .out1({ S4986 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_226_ (
  .in1({ S4986 }),
  .out1({ S4997 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_227_ (
  .in1({ S4975, new_datapath_muxmem_in2_8 }),
  .out1({ S5007 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_228_ (
  .in1({ S5007, S4997 }),
  .out1({ S5018 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_229_ (
  .in1({ new_controller_fib_1, S2985 }),
  .out1({ S5029 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_230_ (
  .in1({ new_controller_fib_2, new_controller_fib_0 }),
  .out1({ S5039 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_231_ (
  .in1({ S5039, new_controller_fib_1 }),
  .out1({ S5050 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_232_ (
  .in1({ S5029, new_controller_fib_2 }),
  .out1({ S5061 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_233_ (
  .in1({ S5050, S3117 }),
  .out1({ S5072 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_234_ (
  .in1({ S5072, S4519 }),
  .out1({ S5082 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_235_ (
  .in1({ S5082 }),
  .out1({ S5093 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_236_ (
  .in1({ S4238, S3969 }),
  .out1({ S5104 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_237_ (
  .in1({ S3892, S3771 }),
  .out1({ S5115 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_238_ (
  .in1({ S3881, S3761 }),
  .out1({ S5125 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_239_ (
  .in1({ S3095, new_controller_opcode_7 }),
  .out1({ S5136 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_240_ (
  .in1({ new_controller_opcode_6, S2592 }),
  .out1({ S5147 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_241_ (
  .in1({ S5147, S4232 }),
  .out1({ S5157 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_242_ (
  .in1({ S5136, S4237 }),
  .out1({ S5168 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_243_ (
  .in1({ S5157, S5115 }),
  .out1({ S5179 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_244_ (
  .in1({ S5179, S5104 }),
  .out1({ S5190 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_245_ (
  .in1({ S3969, S3848 }),
  .out1({ S5200 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_246_ (
  .in1({ S5200, S4570 }),
  .out1({ S5211 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_247_ (
  .in1({ S5211 }),
  .out1({ S5222 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_248_ (
  .in1({ S5222, new_controller_234_B_0 }),
  .out1({ S5232 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_249_ (
  .in1({ S5147, S3914 }),
  .out1({ S5239 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_250_ (
  .in1({ S5136, S3903 }),
  .out1({ S5247 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_251_ (
  .in1({ S3914, S3782 }),
  .out1({ S5255 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_252_ (
  .in1({ S3903, S3793 }),
  .out1({ S5262 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_253_ (
  .in1({ new_controller_opcode_6, S2592 }),
  .out1({ S5271 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_254_ (
  .in1({ S3095, new_controller_opcode_7 }),
  .out1({ S5280 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_255_ (
  .in1({ S5280, S3826 }),
  .out1({ S5290 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_256_ (
  .in1({ S5271, S3815 }),
  .out1({ S5300 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_257_ (
  .in1({ S5290, S5255 }),
  .out1({ S5311 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_258_ (
  .in1({ S5300, S5262 }),
  .out1({ S5322 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_259_ (
  .in1({ S5311, S5247 }),
  .out1({ S5332 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_260_ (
  .in1({ S5322, S3761 }),
  .out1({ S5343 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_261_ (
  .in1({ S5332, S3761 }),
  .out1({ S5354 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_262_ (
  .in1({ S5354 }),
  .out1({ S5365 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_263_ (
  .in1({ S5354, S5232 }),
  .out1({ S5376 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_264_ (
  .in1({ S5376, S5190 }),
  .out1({ S5387 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_265_ (
  .in1({ S5093, S4578 }),
  .out1({ S5398 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_266_ (
  .in1({ S5398, S3969 }),
  .out1({ S5408 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_267_ (
  .in1({ S5408 }),
  .out1({ S5419 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_268_ (
  .in1({ S5408, S5387 }),
  .out1({ S5430 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_269_ (
  .in1({ S5430, new_datapath_instruction_3 }),
  .out1({ S5440 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_270_ (
  .in1({ S3826, S3598 }),
  .out1({ S5451 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_271_ (
  .in1({ S3815, S3587 }),
  .out1({ S5462 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_272_ (
  .in1({ S5280, S4078 }),
  .out1({ S5473 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_273_ (
  .in1({ S5271, S4089 }),
  .out1({ S5483 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_274_ (
  .in1({ S5473, S5451 }),
  .out1({ S5494 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_275_ (
  .in1({ S5483, S5462 }),
  .out1({ S5505 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_276_ (
  .in1({ S5494, S3771 }),
  .out1({ S5515 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_277_ (
  .in1({ S5505, S3761 }),
  .out1({ S5526 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_278_ (
  .in1({ S4563, S3620 }),
  .out1({ S5537 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_279_ (
  .in1({ S4552, S3609 }),
  .out1({ S5547 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_280_ (
  .in1({ S3761, new_controller_opcode_4 }),
  .out1({ S5558 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_281_ (
  .in1({ S5558 }),
  .out1({ S5568 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_282_ (
  .in1({ S4563, S4067 }),
  .out1({ S5579 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_283_ (
  .in1({ S4552, S4056 }),
  .out1({ S5590 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_284_ (
  .in1({ S4563, S4078 }),
  .out1({ S5600 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_285_ (
  .in1({ S4552, S4089 }),
  .out1({ S5611 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_286_ (
  .in1({ S5280, S3914 }),
  .out1({ S5621 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_287_ (
  .in1({ S5271, S3903 }),
  .out1({ S5632 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_288_ (
  .in1({ S5147, S3826 }),
  .out1({ S5642 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_289_ (
  .in1({ S5136, S3815 }),
  .out1({ S5653 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_290_ (
  .in1({ S5642, S5621 }),
  .out1({ S5663 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_291_ (
  .in1({ S5653, S5632 }),
  .out1({ S5673 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_292_ (
  .in1({ S5663, S3771 }),
  .out1({ S5683 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_293_ (
  .in1({ S5673, S3761 }),
  .out1({ S5693 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_294_ (
  .in1({ S5683, S5600 }),
  .out1({ S5702 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_295_ (
  .in1({ S5693, S5611 }),
  .out1({ S5710 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_296_ (
  .in1({ S5710, S5515 }),
  .out1({ S5719 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_297_ (
  .in1({ S5702, S5526 }),
  .out1({ S5729 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_298_ (
  .in1({ S4246, new_controller_opcode_2 }),
  .out1({ S5739 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_299_ (
  .in1({ S5739, S6216 }),
  .out1({ S5749 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_300_ (
  .in1({ S5211, new_controller_234_B_0 }),
  .out1({ S5759 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_301_ (
  .in1({ S5759, S5729 }),
  .out1({ S5770 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_302_ (
  .in1({ S5770, S5749 }),
  .out1({ S5780 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_303_ (
  .in1({ S5780, new_controller_fib_3 }),
  .out1({ S5791 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_304_ (
  .in1({ S5791, S5440 }),
  .out1({ new_datapath_muxrs1_outmux_3 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_305_ (
  .in1({ S5430, new_datapath_instruction_0 }),
  .out1({ S5810 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_306_ (
  .in1({ S5780, new_controller_fib_0 }),
  .out1({ S5821 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_307_ (
  .in1({ S5821, S5810 }),
  .out1({ new_datapath_muxrs1_outmux_0 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_308_ (
  .in1({ new_datapath_muxrs1_outmux_0, new_datapath_muxrs1_outmux_3 }),
  .out1({ S5841 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_309_ (
  .in1({ S5430, new_datapath_instruction_1 }),
  .out1({ S5852 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_310_ (
  .in1({ S5780, new_controller_fib_1 }),
  .out1({ S5862 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_311_ (
  .in1({ S5862, S5852 }),
  .out1({ new_datapath_muxrs1_outmux_1 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_312_ (
  .in1({ S5430, new_datapath_instruction_2 }),
  .out1({ S5882 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_313_ (
  .in1({ S5780, new_controller_fib_2 }),
  .out1({ S5893 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_314_ (
  .in1({ S5893, S5882 }),
  .out1({ new_datapath_muxrs1_outmux_2 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_315_ (
  .in1({ new_datapath_muxrs1_outmux_2, new_datapath_muxrs1_outmux_1 }),
  .out1({ S5902 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_316_ (
  .in1({ S5902, S5841 }),
  .out1({ S5903 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_317_ (
  .in1({ S5903, new_controller_outflag_7 }),
  .out1({ S5904 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_318_ (
  .in1({ S5904 }),
  .out1({ S5905 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_319_ (
  .in1({ S5903, S3226 }),
  .out1({ S5906 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_320_ (
  .in1({ S5906, S5905 }),
  .out1({ S5907 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_321_ (
  .in1({ S5907 }),
  .out1({ new_datapath_addsubunit_in1_7 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_322_ (
  .in1({ new_datapath_addsubunit_in1_7, S4602 }),
  .out1({ S5908 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_323_ (
  .in1({ S5908, S4300 }),
  .out1({ S5909 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_324_ (
  .in1({ S5909, new_datapath_muxmem_in2_7 }),
  .out1({ S5910 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_325_ (
  .in1({ S5910 }),
  .out1({ S5911 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_326_ (
  .in1({ S5909, new_datapath_muxmem_in2_7 }),
  .out1({ S5912 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_327_ (
  .in1({ S5903, new_controller_outflag_6 }),
  .out1({ S5913 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_328_ (
  .in1({ S5913 }),
  .out1({ S5914 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_329_ (
  .in1({ S5903, S3215 }),
  .out1({ S5915 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_330_ (
  .in1({ S5915, S5914 }),
  .out1({ S5916 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_331_ (
  .in1({ S5916 }),
  .out1({ new_datapath_addsubunit_in1_6 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_332_ (
  .in1({ new_datapath_addsubunit_in1_6, S4602 }),
  .out1({ S5917 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_333_ (
  .in1({ S5917, S4300 }),
  .out1({ S5918 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_334_ (
  .in1({ S5918, new_datapath_muxmem_in2_6 }),
  .out1({ S5919 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_335_ (
  .in1({ S5919 }),
  .out1({ S5920 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_336_ (
  .in1({ S5918, new_datapath_muxmem_in2_6 }),
  .out1({ S5921 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_337_ (
  .in1({ S5921, S5920 }),
  .out1({ S5922 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_338_ (
  .in1({ S5903, new_controller_407_B_2 }),
  .out1({ S5923 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_339_ (
  .in1({ S5923 }),
  .out1({ S5924 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_340_ (
  .in1({ S5903, S3204 }),
  .out1({ S5925 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_341_ (
  .in1({ S5925, S5924 }),
  .out1({ S5926 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_342_ (
  .in1({ S5926 }),
  .out1({ new_datapath_addsubunit_in1_5 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_343_ (
  .in1({ new_datapath_addsubunit_in1_5, S4602 }),
  .out1({ S5927 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_344_ (
  .in1({ S5927, S4300 }),
  .out1({ S5928 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_345_ (
  .in1({ S5928, new_datapath_muxmem_in2_5 }),
  .out1({ S5929 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_346_ (
  .in1({ S5929 }),
  .out1({ S5930 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_347_ (
  .in1({ S5928, new_datapath_muxmem_in2_5 }),
  .out1({ S5931 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_348_ (
  .in1({ S4289, new_controller_fib_4 }),
  .out1({ S5932 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_349_ (
  .in1({ S5903, new_controller_407_B_0 }),
  .out1({ S5933 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_350_ (
  .in1({ S5933 }),
  .out1({ S5934 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_351_ (
  .in1({ S5903, S3193 }),
  .out1({ S5935 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_352_ (
  .in1({ S5935, S5934 }),
  .out1({ S5936 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_353_ (
  .in1({ S5936 }),
  .out1({ new_datapath_addsubunit_in1_4 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_354_ (
  .in1({ new_datapath_addsubunit_in1_4, S4602 }),
  .out1({ S5937 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_355_ (
  .in1({ S5937, S5932 }),
  .out1({ S5938 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_356_ (
  .in1({ S5938, new_datapath_muxmem_in2_4 }),
  .out1({ S5939 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_357_ (
  .in1({ S5939 }),
  .out1({ S5940 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_358_ (
  .in1({ S5938, new_datapath_muxmem_in2_4 }),
  .out1({ S5941 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_359_ (
  .in1({ S5941, S5940 }),
  .out1({ S5942 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_360_ (
  .in1({ S4289, new_controller_fib_3 }),
  .out1({ S5943 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_361_ (
  .in1({ S5903, new_controller_outflag_3 }),
  .out1({ S5944 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_362_ (
  .in1({ S5944 }),
  .out1({ S5945 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_363_ (
  .in1({ S5903, S3182 }),
  .out1({ S5946 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_364_ (
  .in1({ S5946, S5945 }),
  .out1({ S5947 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_365_ (
  .in1({ S5947 }),
  .out1({ new_datapath_addsubunit_in1_3 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_366_ (
  .in1({ new_datapath_addsubunit_in1_3, S4602 }),
  .out1({ S5948 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_367_ (
  .in1({ S5948, S5943 }),
  .out1({ S5949 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_368_ (
  .in1({ S5949, new_datapath_muxmem_in2_3 }),
  .out1({ S5950 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_369_ (
  .in1({ S5950 }),
  .out1({ S5951 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_370_ (
  .in1({ S5949, new_datapath_muxmem_in2_3 }),
  .out1({ S5952 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_371_ (
  .in1({ S4289, new_controller_fib_2 }),
  .out1({ S5953 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_372_ (
  .in1({ S5903, new_controller_outflag_2 }),
  .out1({ S5954 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_373_ (
  .in1({ S5954 }),
  .out1({ S5955 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_374_ (
  .in1({ S5903, S3171 }),
  .out1({ S5956 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_375_ (
  .in1({ S5956, S5955 }),
  .out1({ S5957 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_376_ (
  .in1({ S5957 }),
  .out1({ new_datapath_addsubunit_in1_2 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_377_ (
  .in1({ new_datapath_addsubunit_in1_2, S4602 }),
  .out1({ S5958 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_378_ (
  .in1({ S5958, S5953 }),
  .out1({ S5959 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_379_ (
  .in1({ S5959, new_datapath_muxmem_in2_2 }),
  .out1({ S5960 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_380_ (
  .in1({ S5960 }),
  .out1({ S5961 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_381_ (
  .in1({ S4289, new_controller_fib_1 }),
  .out1({ S5962 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_382_ (
  .in1({ S5903, new_controller_outflag_1 }),
  .out1({ S5963 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_383_ (
  .in1({ S5963 }),
  .out1({ S5964 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_384_ (
  .in1({ S5903, S3160 }),
  .out1({ S5965 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_385_ (
  .in1({ S5965, S5964 }),
  .out1({ S5966 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_386_ (
  .in1({ S5966 }),
  .out1({ new_datapath_addsubunit_in1_1 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_387_ (
  .in1({ new_datapath_addsubunit_in1_1, S4602 }),
  .out1({ S5967 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_388_ (
  .in1({ S5967, S5962 }),
  .out1({ S5968 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_389_ (
  .in1({ S5968, new_datapath_muxmem_in2_1 }),
  .out1({ S5969 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_390_ (
  .in1({ S5969 }),
  .out1({ S5970 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_391_ (
  .in1({ S4289, new_controller_fib_0 }),
  .out1({ S5971 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_392_ (
  .in1({ S5903, new_controller_outflag_0 }),
  .out1({ S5972 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_393_ (
  .in1({ S5972 }),
  .out1({ S5973 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_394_ (
  .in1({ S5903, S3150 }),
  .out1({ S5974 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_395_ (
  .in1({ S5974, S5973 }),
  .out1({ S5975 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_396_ (
  .in1({ S5975 }),
  .out1({ new_datapath_addsubunit_in1_0 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_397_ (
  .in1({ new_datapath_addsubunit_in1_0, S4602 }),
  .out1({ S5976 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_398_ (
  .in1({ S5976, S5971 }),
  .out1({ S5977 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_399_ (
  .in1({ S5977 }),
  .out1({ S5978 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_400_ (
  .in1({ S5978, S2625 }),
  .out1({ S5979 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_401_ (
  .in1({ S5968, new_datapath_muxmem_in2_1 }),
  .out1({ S5980 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_402_ (
  .in1({ S5980, S5970 }),
  .out1({ S5981 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_403_ (
  .in1({ S5981, S5979 }),
  .out1({ S5982 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_404_ (
  .in1({ S5982, S5969 }),
  .out1({ S5983 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_405_ (
  .in1({ S5959, new_datapath_muxmem_in2_2 }),
  .out1({ S5984 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_406_ (
  .in1({ S5984, S5961 }),
  .out1({ S5985 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_407_ (
  .in1({ S5985, S5983 }),
  .out1({ S5986 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_408_ (
  .in1({ S5986, S5960 }),
  .out1({ S5987 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_409_ (
  .in1({ S5987, S5951 }),
  .out1({ S5988 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_410_ (
  .in1({ S5988, S5952 }),
  .out1({ S5989 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_411_ (
  .in1({ S5989, S5942 }),
  .out1({ S5990 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_412_ (
  .in1({ S5990, S5939 }),
  .out1({ S5991 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_413_ (
  .in1({ S5991, S5930 }),
  .out1({ S5992 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_414_ (
  .in1({ S5992, S5931 }),
  .out1({ S5993 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_415_ (
  .in1({ S5993, S5922 }),
  .out1({ S5994 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_416_ (
  .in1({ S5994, S5919 }),
  .out1({ S5995 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_417_ (
  .in1({ S5995, S5911 }),
  .out1({ S5996 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_418_ (
  .in1({ S5996, S5912 }),
  .out1({ S5997 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_419_ (
  .in1({ S5997, S5018 }),
  .out1({ S5998 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_420_ (
  .in1({ S5998, S4986 }),
  .out1({ S5999 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_421_ (
  .in1({ S5999, S4943 }),
  .out1({ S6000 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_422_ (
  .in1({ S6000, S4954 }),
  .out1({ S6001 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_423_ (
  .in1({ S6001, S4900 }),
  .out1({ S6002 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_424_ (
  .in1({ S6002, S4868 }),
  .out1({ S6003 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_425_ (
  .in1({ S6003, S4836 }),
  .out1({ S6004 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_426_ (
  .in1({ S6004, S4825 }),
  .out1({ S6005 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_427_ (
  .in1({ S6005, S4783 }),
  .out1({ S6006 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_428_ (
  .in1({ S6006, S4750 }),
  .out1({ S6007 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_429_ (
  .in1({ S6007, S4708 }),
  .out1({ S6008 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_430_ (
  .in1({ S6008, S4718 }),
  .out1({ S6009 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_431_ (
  .in1({ S6009, S4665 }),
  .out1({ S6010 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_432_ (
  .in1({ S6010, S4632 }),
  .out1({ S6011 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_433_ (
  .in1({ S4602, new_datapath_addsubunit_in1_15 }),
  .out1({ S6012 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_434_ (
  .in1({ S6012, S4300 }),
  .out1({ S6013 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_435_ (
  .in1({ S6013, new_datapath_muxmem_in2_15 }),
  .out1({ S6014 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_436_ (
  .in1({ S6014 }),
  .out1({ S6015 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_437_ (
  .in1({ S6013, new_datapath_muxmem_in2_15 }),
  .out1({ S6016 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_438_ (
  .in1({ S6016, S6015 }),
  .out1({ S6017 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_439_ (
  .in1({ S6017, S6011 }),
  .out1({ S6018 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_440_ (
  .in1({ S5082, S4586 }),
  .out1({ S6019 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_441_ (
  .in1({ S6019 }),
  .out1({ S6020 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_442_ (
  .in1({ S6020, S4254 }),
  .out1({ S6021 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_443_ (
  .in1({ S6017, S6011 }),
  .out1({ S6022 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_444_ (
  .in1({ S6021, S6018 }),
  .out1({ S6023 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_445_ (
  .in1({ S6023, S6022 }),
  .out1({ S6024 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_446_ (
  .in1({ S4399, new_controller_407_B_0 }),
  .out1({ S6025 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_447_ (
  .in1({ S6025, S4443 }),
  .out1({ S6026 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_448_ (
  .in1({ S6026, S4344 }),
  .out1({ S6027 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_449_ (
  .in1({ S4487, new_controller_407_B_0 }),
  .out1({ S6028 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_450_ (
  .in1({ S4421, S4344 }),
  .out1({ S6029 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_451_ (
  .in1({ S6029, S2996 }),
  .out1({ S6030 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_452_ (
  .in1({ S6030, S6028 }),
  .out1({ S6031 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_453_ (
  .in1({ S5061, S3117 }),
  .out1({ S6032 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_454_ (
  .in1({ S4355, S4322 }),
  .out1({ S6033 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_455_ (
  .in1({ S6033, S3969 }),
  .out1({ S6034 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_456_ (
  .in1({ S6034, S6032 }),
  .out1({ S6035 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_457_ (
  .in1({ S6035, S6031 }),
  .out1({ S6036 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_458_ (
  .in1({ S6036, S6027 }),
  .out1({ S6037 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_459_ (
  .in1({ S6037, S3958 }),
  .out1({ S6038 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_460_ (
  .in1({ S6038, S3936 }),
  .out1({ S6039 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_461_ (
  .in1({ S6039, S3771 }),
  .out1({ S6040 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_462_ (
  .in1({ S4155, S3719 }),
  .out1({ S6041 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_463_ (
  .in1({ S6041, S6040 }),
  .out1({ S6042 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_464_ (
  .in1({ S2636, S2625 }),
  .out1({ S6043 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_465_ (
  .in1({ new_datapath_muxmem_in2_1, new_datapath_muxmem_in2_0 }),
  .out1({ S6044 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_466_ (
  .in1({ S6044, S2647 }),
  .out1({ S6045 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_467_ (
  .in1({ S6043, new_datapath_muxmem_in2_2 }),
  .out1({ S6046 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_468_ (
  .in1({ S6046, S2658 }),
  .out1({ S6047 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_469_ (
  .in1({ S6045, new_datapath_muxmem_in2_3 }),
  .out1({ S6048 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_470_ (
  .in1({ S6047, new_datapath_muxmem_in2_4 }),
  .out1({ S6049 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_471_ (
  .in1({ S6049 }),
  .out1({ S6050 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_472_ (
  .in1({ S6050, new_datapath_muxmem_in2_5 }),
  .out1({ S6051 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_473_ (
  .in1({ S6051 }),
  .out1({ S6052 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_474_ (
  .in1({ S6052, new_datapath_muxmem_in2_6 }),
  .out1({ S6053 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_475_ (
  .in1({ S6053 }),
  .out1({ S6054 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_476_ (
  .in1({ S6054, new_datapath_muxmem_in2_7 }),
  .out1({ S6055 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_477_ (
  .in1({ S6055 }),
  .out1({ S6056 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_478_ (
  .in1({ S6055, S2712 }),
  .out1({ S6057 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_479_ (
  .in1({ S6056, new_datapath_muxmem_in2_8 }),
  .out1({ S6058 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_480_ (
  .in1({ S6058, S2723 }),
  .out1({ S6059 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_481_ (
  .in1({ S6057, new_datapath_muxmem_in2_9 }),
  .out1({ S6060 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_482_ (
  .in1({ S6060, S2734 }),
  .out1({ S6061 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_483_ (
  .in1({ S6059, new_datapath_muxmem_in2_10 }),
  .out1({ S6062 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_484_ (
  .in1({ S6061, new_datapath_muxmem_in2_11 }),
  .out1({ S6063 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_485_ (
  .in1({ S6063 }),
  .out1({ S6064 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_486_ (
  .in1({ S6064, new_datapath_muxmem_in2_12 }),
  .out1({ S6065 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_487_ (
  .in1({ S6065 }),
  .out1({ S6066 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_488_ (
  .in1({ S6065, S2767 }),
  .out1({ S6067 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_489_ (
  .in1({ S6066, new_datapath_muxmem_in2_13 }),
  .out1({ S6068 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_490_ (
  .in1({ S6067, new_datapath_muxmem_in2_14 }),
  .out1({ S6069 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_491_ (
  .in1({ S6069 }),
  .out1({ S6070 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_492_ (
  .in1({ S6069, new_datapath_muxmem_in2_15 }),
  .out1({ S6071 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_493_ (
  .in1({ S6069, new_datapath_muxmem_in2_15 }),
  .out1({ S6072 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_494_ (
  .in1({ S6072 }),
  .out1({ S6073 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_495_ (
  .in1({ S6073, S6071 }),
  .out1({ S6074 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_496_ (
  .in1({ S6074 }),
  .out1({ S6075 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_497_ (
  .in1({ S6075, S6042 }),
  .out1({ S6076 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_498_ (
  .in1({ S5072, new_controller_234_B_0 }),
  .out1({ S6077 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_499_ (
  .in1({ S6077 }),
  .out1({ S6078 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_500_ (
  .in1({ S6078, S5408 }),
  .out1({ S6079 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_501_ (
  .in1({ S6077, S5419 }),
  .out1({ S6080 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_502_ (
  .in1({ S6079, S6076 }),
  .out1({ S6081 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_503_ (
  .in1({ S6081, S6024 }),
  .out1({ S6082 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_504_ (
  .in1({ S6080, new_datapath_addsubunit_in1_15 }),
  .out1({ S6083 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_505_ (
  .in1({ S6083, S4210 }),
  .out1({ S6084 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_506_ (
  .in1({ S6084, S6082 }),
  .out1({ S6085 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_507_ (
  .in1({ S6085, S4221 }),
  .out1({ S0 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_508_ (
  .in1({ S4133, new_controller_pstate_0 }),
  .out1({ S6086 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_509_ (
  .in1({ S6086, S2581 }),
  .out1({ S1 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_510_ (
  .in1({ S3139, S3128 }),
  .out1({ S6087 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_511_ (
  .in1({ S6087 }),
  .out1({ new_controller_1133_S_0 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_512_ (
  .in1({ new_controller_1133_S_0, new_datapath_databusin_15 }),
  .out1({ S6088 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_513_ (
  .in1({ S6087, new_controller_opcode_7 }),
  .out1({ S6089 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_514_ (
  .in1({ S6089, S6088 }),
  .out1({ S2 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_515_ (
  .in1({ S4246, new_controller_opcode_3 }),
  .out1({ S6090 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_516_ (
  .in1({ S4238, S3062 }),
  .out1({ S6091 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_517_ (
  .in1({ S6091, new_datapath_adr_outreg_15 }),
  .out1({ S6092 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_518_ (
  .in1({ S6090, S6013 }),
  .out1({ S6093 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_519_ (
  .in1({ S6093, S6092 }),
  .out1({ S4 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_520_ (
  .in1({ S4210, new_datapath_muxmem_in2_0 }),
  .out1({ S6094 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_521_ (
  .in1({ S5978, S2625 }),
  .out1({ S6095 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_522_ (
  .in1({ S6021, S5979 }),
  .out1({ S6096 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_523_ (
  .in1({ S6096, S6095 }),
  .out1({ S6097 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_524_ (
  .in1({ S6042, new_datapath_muxmem_in2_0 }),
  .out1({ S6098 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_525_ (
  .in1({ S6098, S6079 }),
  .out1({ S6099 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_526_ (
  .in1({ S6099, S6097 }),
  .out1({ S6100 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_527_ (
  .in1({ S6080, new_datapath_addsubunit_in1_0 }),
  .out1({ S6101 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_528_ (
  .in1({ S6101, S4210 }),
  .out1({ S6102 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_529_ (
  .in1({ S6102, S6100 }),
  .out1({ S6103 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_530_ (
  .in1({ S6103, S6094 }),
  .out1({ S5 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_531_ (
  .in1({ S4210, new_datapath_muxmem_in2_1 }),
  .out1({ S6104 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_532_ (
  .in1({ S5981, S5979 }),
  .out1({ S6105 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_533_ (
  .in1({ S6105, S6021 }),
  .out1({ S6106 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_534_ (
  .in1({ S6106, S5982 }),
  .out1({ S6107 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_535_ (
  .in1({ new_datapath_muxmem_in2_1, new_datapath_muxmem_in2_0 }),
  .out1({ S6108 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_536_ (
  .in1({ S6108 }),
  .out1({ S6109 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_537_ (
  .in1({ S6108, S6043 }),
  .out1({ S6110 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_538_ (
  .in1({ S6109, S6044 }),
  .out1({ S6111 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_539_ (
  .in1({ S6111, S6042 }),
  .out1({ S6112 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_540_ (
  .in1({ S6112, S6079 }),
  .out1({ S6113 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_541_ (
  .in1({ S6113, S6107 }),
  .out1({ S6114 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_542_ (
  .in1({ S6080, new_datapath_addsubunit_in1_1 }),
  .out1({ S6115 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_543_ (
  .in1({ S6115, S4210 }),
  .out1({ S6116 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_544_ (
  .in1({ S6116, S6114 }),
  .out1({ S6117 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_545_ (
  .in1({ S6117, S6104 }),
  .out1({ S6 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_546_ (
  .in1({ S4210, new_datapath_muxmem_in2_2 }),
  .out1({ S6118 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_547_ (
  .in1({ S5985, S5983 }),
  .out1({ S6119 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_548_ (
  .in1({ S6119, S6021 }),
  .out1({ S6120 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_549_ (
  .in1({ S6120, S5986 }),
  .out1({ S6121 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_550_ (
  .in1({ S6043, new_datapath_muxmem_in2_2 }),
  .out1({ S6122 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_551_ (
  .in1({ S6044, S2647 }),
  .out1({ S6123 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_552_ (
  .in1({ S6122, S6045 }),
  .out1({ S6124 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_553_ (
  .in1({ S6123, S6046 }),
  .out1({ S6125 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_554_ (
  .in1({ S6125, S6042 }),
  .out1({ S6126 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_555_ (
  .in1({ S6126, S6079 }),
  .out1({ S6127 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_556_ (
  .in1({ S6127, S6121 }),
  .out1({ S6128 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_557_ (
  .in1({ S6080, new_datapath_addsubunit_in1_2 }),
  .out1({ S6129 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_558_ (
  .in1({ S6129, S4210 }),
  .out1({ S6130 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_559_ (
  .in1({ S6130, S6128 }),
  .out1({ S6131 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_560_ (
  .in1({ S6131, S6118 }),
  .out1({ S7 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_561_ (
  .in1({ S4210, new_datapath_muxmem_in2_3 }),
  .out1({ S6132 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_562_ (
  .in1({ S5952, S5951 }),
  .out1({ S6133 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_563_ (
  .in1({ S6133, S5987 }),
  .out1({ S6134 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_564_ (
  .in1({ S6133, S5987 }),
  .out1({ S6135 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_565_ (
  .in1({ S6135, S6021 }),
  .out1({ S6136 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_566_ (
  .in1({ S6136, S6134 }),
  .out1({ S6137 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_567_ (
  .in1({ S6045, new_datapath_muxmem_in2_3 }),
  .out1({ S6138 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_568_ (
  .in1({ S6046, S2658 }),
  .out1({ S6139 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_569_ (
  .in1({ S6138, S6047 }),
  .out1({ S6140 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_570_ (
  .in1({ S6139, S6048 }),
  .out1({ S6141 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_571_ (
  .in1({ S6141, S6042 }),
  .out1({ S6142 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_572_ (
  .in1({ S6142, S6079 }),
  .out1({ S6143 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_573_ (
  .in1({ S6143, S6137 }),
  .out1({ S6144 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_574_ (
  .in1({ S6080, new_datapath_addsubunit_in1_3 }),
  .out1({ S6145 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_575_ (
  .in1({ S6145, S4210 }),
  .out1({ S6146 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_576_ (
  .in1({ S6146, S6144 }),
  .out1({ S6147 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_577_ (
  .in1({ S6147, S6132 }),
  .out1({ S8 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_578_ (
  .in1({ S4210, new_datapath_muxmem_in2_4 }),
  .out1({ S6148 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_579_ (
  .in1({ S5989, S5942 }),
  .out1({ S6149 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_580_ (
  .in1({ S6149, S6021 }),
  .out1({ S6150 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_581_ (
  .in1({ S6150, S5990 }),
  .out1({ S6151 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_582_ (
  .in1({ S6048, S2669 }),
  .out1({ S6152 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_583_ (
  .in1({ S6152, S6049 }),
  .out1({ S6153 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_584_ (
  .in1({ S6153, S6042 }),
  .out1({ S6154 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_585_ (
  .in1({ S6154, S6079 }),
  .out1({ S6155 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_586_ (
  .in1({ S6155, S6151 }),
  .out1({ S6156 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_587_ (
  .in1({ S6080, new_datapath_addsubunit_in1_4 }),
  .out1({ S6157 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_588_ (
  .in1({ S6157, S4210 }),
  .out1({ S6158 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_589_ (
  .in1({ S6158, S6156 }),
  .out1({ S6159 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_590_ (
  .in1({ S6159, S6148 }),
  .out1({ S9 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_591_ (
  .in1({ S4210, new_datapath_muxmem_in2_5 }),
  .out1({ S6160 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_592_ (
  .in1({ S5931, S5930 }),
  .out1({ S6161 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_593_ (
  .in1({ S6161, S5991 }),
  .out1({ S6162 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_594_ (
  .in1({ S6161, S5991 }),
  .out1({ S6163 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_595_ (
  .in1({ S6163, S6021 }),
  .out1({ S6164 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_596_ (
  .in1({ S6164, S6162 }),
  .out1({ S6165 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_597_ (
  .in1({ S6049, S2680 }),
  .out1({ S6166 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_598_ (
  .in1({ S6166, S6051 }),
  .out1({ S6167 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_599_ (
  .in1({ S6167, S6042 }),
  .out1({ S6168 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_600_ (
  .in1({ S6168, S6079 }),
  .out1({ S6169 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_601_ (
  .in1({ S6169, S6165 }),
  .out1({ S6170 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_602_ (
  .in1({ S6080, new_datapath_addsubunit_in1_5 }),
  .out1({ S6171 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_603_ (
  .in1({ S6171, S4210 }),
  .out1({ S6172 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_604_ (
  .in1({ S6172, S6170 }),
  .out1({ S6173 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_605_ (
  .in1({ S6173, S6160 }),
  .out1({ S10 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_606_ (
  .in1({ S4210, new_datapath_muxmem_in2_6 }),
  .out1({ S6174 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_607_ (
  .in1({ S5993, S5922 }),
  .out1({ S6175 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_608_ (
  .in1({ S6175, S6021 }),
  .out1({ S6176 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_609_ (
  .in1({ S6176, S5994 }),
  .out1({ S6177 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_610_ (
  .in1({ S6051, S2690 }),
  .out1({ S6178 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_611_ (
  .in1({ S6178, S6053 }),
  .out1({ S6179 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_612_ (
  .in1({ S6179, S6042 }),
  .out1({ S6180 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_613_ (
  .in1({ S6180, S6079 }),
  .out1({ S6181 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_614_ (
  .in1({ S6181, S6177 }),
  .out1({ S6182 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_615_ (
  .in1({ S6080, new_datapath_addsubunit_in1_6 }),
  .out1({ S6183 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_616_ (
  .in1({ S6183, S4210 }),
  .out1({ S6184 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_617_ (
  .in1({ S6184, S6182 }),
  .out1({ S6185 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_618_ (
  .in1({ S6185, S6174 }),
  .out1({ S11 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_619_ (
  .in1({ S4210, new_datapath_muxmem_in2_7 }),
  .out1({ S6186 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_620_ (
  .in1({ S5912, S5911 }),
  .out1({ S6187 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_621_ (
  .in1({ S6187, S5995 }),
  .out1({ S6188 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_622_ (
  .in1({ S6187, S5995 }),
  .out1({ S6189 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_623_ (
  .in1({ S6189, S6021 }),
  .out1({ S6190 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_624_ (
  .in1({ S6190, S6188 }),
  .out1({ S6191 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_625_ (
  .in1({ S6053, S2701 }),
  .out1({ S6192 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_626_ (
  .in1({ S6192, S6055 }),
  .out1({ S6193 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_627_ (
  .in1({ S6193, S6042 }),
  .out1({ S6194 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_628_ (
  .in1({ S6194, S6079 }),
  .out1({ S6195 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_629_ (
  .in1({ S6195, S6191 }),
  .out1({ S6196 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_630_ (
  .in1({ S6080, new_datapath_addsubunit_in1_7 }),
  .out1({ S6197 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_631_ (
  .in1({ S6197, S4210 }),
  .out1({ S6198 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_632_ (
  .in1({ S6198, S6196 }),
  .out1({ S6199 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_633_ (
  .in1({ S6199, S6186 }),
  .out1({ S12 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_634_ (
  .in1({ S4210, new_datapath_muxmem_in2_8 }),
  .out1({ S6200 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_635_ (
  .in1({ S5997, S5018 }),
  .out1({ S6201 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_636_ (
  .in1({ S6201, S6021 }),
  .out1({ S6202 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_637_ (
  .in1({ S6202, S5998 }),
  .out1({ S6203 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_638_ (
  .in1({ S6055, S2712 }),
  .out1({ S6204 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_639_ (
  .in1({ S6204, S6058 }),
  .out1({ S6205 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_640_ (
  .in1({ S6205, S6042 }),
  .out1({ S6206 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_641_ (
  .in1({ S6206, S6079 }),
  .out1({ S6207 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_642_ (
  .in1({ S6207, S6203 }),
  .out1({ S6208 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_643_ (
  .in1({ S6080, new_datapath_addsubunit_in1_8 }),
  .out1({ S6209 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_644_ (
  .in1({ S6209, S4210 }),
  .out1({ S6210 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_645_ (
  .in1({ S6210, S6208 }),
  .out1({ S6211 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_646_ (
  .in1({ S6211, S6200 }),
  .out1({ S13 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_647_ (
  .in1({ S4210, new_datapath_muxmem_in2_9 }),
  .out1({ S6212 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_648_ (
  .in1({ S4954, S4943 }),
  .out1({ S6213 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_649_ (
  .in1({ S6213, S5999 }),
  .out1({ S6214 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_650_ (
  .in1({ S6213, S5999 }),
  .out1({ S88 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_651_ (
  .in1({ S88, S6021 }),
  .out1({ S89 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_652_ (
  .in1({ S89, S6214 }),
  .out1({ S90 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_653_ (
  .in1({ S6057, new_datapath_muxmem_in2_9 }),
  .out1({ S91 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_654_ (
  .in1({ S6058, S2723 }),
  .out1({ S92 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_655_ (
  .in1({ S91, S6059 }),
  .out1({ S93 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_656_ (
  .in1({ S92, S6060 }),
  .out1({ S94 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_657_ (
  .in1({ S94, S6042 }),
  .out1({ S95 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_658_ (
  .in1({ S95, S6079 }),
  .out1({ S96 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_659_ (
  .in1({ S96, S90 }),
  .out1({ S97 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_660_ (
  .in1({ S6080, new_datapath_addsubunit_in1_9 }),
  .out1({ S98 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_661_ (
  .in1({ S98, S4210 }),
  .out1({ S99 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_662_ (
  .in1({ S99, S97 }),
  .out1({ S100 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_663_ (
  .in1({ S100, S6212 }),
  .out1({ S14 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_664_ (
  .in1({ S4210, new_datapath_muxmem_in2_10 }),
  .out1({ S101 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_665_ (
  .in1({ S6001, S4900 }),
  .out1({ S102 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_666_ (
  .in1({ S102, S6021 }),
  .out1({ S103 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_667_ (
  .in1({ S103, S6002 }),
  .out1({ S104 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_668_ (
  .in1({ S6059, new_datapath_muxmem_in2_10 }),
  .out1({ S105 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_669_ (
  .in1({ S6060, S2734 }),
  .out1({ S106 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_670_ (
  .in1({ S105, S6061 }),
  .out1({ S107 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_671_ (
  .in1({ S106, S6062 }),
  .out1({ S108 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_672_ (
  .in1({ S108, S6042 }),
  .out1({ S109 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_673_ (
  .in1({ S109, S6079 }),
  .out1({ S110 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_674_ (
  .in1({ S110, S104 }),
  .out1({ S111 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_675_ (
  .in1({ S6080, new_datapath_addsubunit_in1_10 }),
  .out1({ S112 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_676_ (
  .in1({ S112, S4210 }),
  .out1({ S113 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_677_ (
  .in1({ S113, S111 }),
  .out1({ S114 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_678_ (
  .in1({ S114, S101 }),
  .out1({ S15 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_679_ (
  .in1({ S4210, new_datapath_muxmem_in2_11 }),
  .out1({ S115 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_680_ (
  .in1({ S4836, S4825 }),
  .out1({ S116 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_681_ (
  .in1({ S116, S6003 }),
  .out1({ S117 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_682_ (
  .in1({ S116, S6003 }),
  .out1({ S118 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_683_ (
  .in1({ S118, S6021 }),
  .out1({ S119 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_684_ (
  .in1({ S119, S117 }),
  .out1({ S120 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_685_ (
  .in1({ S6062, S2745 }),
  .out1({ S121 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_686_ (
  .in1({ S121, S6063 }),
  .out1({ S122 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_687_ (
  .in1({ S122, S6042 }),
  .out1({ S123 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_688_ (
  .in1({ S123, S6079 }),
  .out1({ S124 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_689_ (
  .in1({ S124, S120 }),
  .out1({ S125 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_690_ (
  .in1({ S6080, new_datapath_addsubunit_in1_11 }),
  .out1({ S126 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_691_ (
  .in1({ S126, S4210 }),
  .out1({ S127 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_692_ (
  .in1({ S127, S125 }),
  .out1({ S128 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_693_ (
  .in1({ S128, S115 }),
  .out1({ S16 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_694_ (
  .in1({ S4210, new_datapath_muxmem_in2_12 }),
  .out1({ S129 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_695_ (
  .in1({ S6005, S4783 }),
  .out1({ S130 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_696_ (
  .in1({ S130, S6021 }),
  .out1({ S131 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_697_ (
  .in1({ S131, S6006 }),
  .out1({ S132 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_698_ (
  .in1({ S6063, S2756 }),
  .out1({ S133 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_699_ (
  .in1({ S133, S6065 }),
  .out1({ S134 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_700_ (
  .in1({ S134, S6042 }),
  .out1({ S135 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_701_ (
  .in1({ S135, S6079 }),
  .out1({ S136 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_702_ (
  .in1({ S136, S132 }),
  .out1({ S137 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_703_ (
  .in1({ S6080, new_datapath_addsubunit_in1_12 }),
  .out1({ S138 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_704_ (
  .in1({ S138, S4210 }),
  .out1({ S139 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_705_ (
  .in1({ S139, S137 }),
  .out1({ S140 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_706_ (
  .in1({ S140, S129 }),
  .out1({ S17 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_707_ (
  .in1({ S4210, new_datapath_muxmem_in2_13 }),
  .out1({ S141 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_708_ (
  .in1({ S4718, S4708 }),
  .out1({ S142 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_709_ (
  .in1({ S142, S6007 }),
  .out1({ S143 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_710_ (
  .in1({ S142, S6007 }),
  .out1({ S144 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_711_ (
  .in1({ S144, S6021 }),
  .out1({ S145 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_712_ (
  .in1({ S145, S143 }),
  .out1({ S146 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_713_ (
  .in1({ S6065, S2767 }),
  .out1({ S147 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_714_ (
  .in1({ S147, S6068 }),
  .out1({ S148 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_715_ (
  .in1({ S148, S6042 }),
  .out1({ S149 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_716_ (
  .in1({ S149, S6079 }),
  .out1({ S150 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_717_ (
  .in1({ S150, S146 }),
  .out1({ S151 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_718_ (
  .in1({ S6080, new_datapath_addsubunit_in1_13 }),
  .out1({ S152 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_719_ (
  .in1({ S152, S4210 }),
  .out1({ S153 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_720_ (
  .in1({ S153, S151 }),
  .out1({ S154 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_721_ (
  .in1({ S154, S141 }),
  .out1({ S18 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_722_ (
  .in1({ S4210, new_datapath_muxmem_in2_14 }),
  .out1({ S155 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_723_ (
  .in1({ S6009, S4665 }),
  .out1({ S156 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_724_ (
  .in1({ S156, S6021 }),
  .out1({ S157 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_725_ (
  .in1({ S157, S6010 }),
  .out1({ S158 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_726_ (
  .in1({ S6067, new_datapath_muxmem_in2_14 }),
  .out1({ S159 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_727_ (
  .in1({ S6068, S2778 }),
  .out1({ S160 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_728_ (
  .in1({ S159, S6070 }),
  .out1({ S161 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_729_ (
  .in1({ S160, S6069 }),
  .out1({ S162 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_730_ (
  .in1({ S162, S6042 }),
  .out1({ S163 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_731_ (
  .in1({ S163, S6079 }),
  .out1({ S164 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_732_ (
  .in1({ S164, S158 }),
  .out1({ S165 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_733_ (
  .in1({ S6080, new_datapath_addsubunit_in1_14 }),
  .out1({ S166 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_734_ (
  .in1({ S166, S4210 }),
  .out1({ S167 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_735_ (
  .in1({ S167, S165 }),
  .out1({ S168 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_736_ (
  .in1({ S168, S155 }),
  .out1({ S19 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_737_ (
  .in1({ S5719, S3062 }),
  .out1({ S169 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_738_ (
  .in1({ new_controller_opcode_2, new_controller_234_B_0 }),
  .out1({ S170 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_739_ (
  .in1({ S4578, new_controller_opcode_3 }),
  .out1({ S171 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_740_ (
  .in1({ S171 }),
  .out1({ S172 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_741_ (
  .in1({ new_controller_opcode_3, new_controller_opcode_2 }),
  .out1({ S173 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_742_ (
  .in1({ S173, S4570 }),
  .out1({ S174 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_743_ (
  .in1({ S174, new_controller_234_B_0 }),
  .out1({ S175 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_744_ (
  .in1({ S175 }),
  .out1({ S176 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_745_ (
  .in1({ S175, new_datapath_instruction_3 }),
  .out1({ S177 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_746_ (
  .in1({ S177 }),
  .out1({ S178 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_747_ (
  .in1({ S178, S169 }),
  .out1({ S179 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_748_ (
  .in1({ S179 }),
  .out1({ new_datapath_muxrs2_outmux_3 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_749_ (
  .in1({ S5719, S3029 }),
  .out1({ S180 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_750_ (
  .in1({ S175, new_datapath_instruction_0 }),
  .out1({ S181 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_751_ (
  .in1({ S181 }),
  .out1({ S182 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_752_ (
  .in1({ S182, S180 }),
  .out1({ S183 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_753_ (
  .in1({ S183 }),
  .out1({ new_datapath_muxrs2_outmux_0 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_754_ (
  .in1({ S183, S179 }),
  .out1({ S184 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_755_ (
  .in1({ new_datapath_muxrs2_outmux_0, new_datapath_muxrs2_outmux_3 }),
  .out1({ S185 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_756_ (
  .in1({ S5719, S3040 }),
  .out1({ S186 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_757_ (
  .in1({ S175, new_datapath_instruction_1 }),
  .out1({ S187 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_758_ (
  .in1({ S187 }),
  .out1({ S188 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_759_ (
  .in1({ S188, S186 }),
  .out1({ S189 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_760_ (
  .in1({ S189 }),
  .out1({ new_datapath_muxrs2_outmux_1 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_761_ (
  .in1({ S5719, S3051 }),
  .out1({ S190 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_762_ (
  .in1({ S175, new_datapath_instruction_2 }),
  .out1({ S191 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_763_ (
  .in1({ S191 }),
  .out1({ S192 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_764_ (
  .in1({ S192, S190 }),
  .out1({ S193 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_765_ (
  .in1({ S193 }),
  .out1({ new_datapath_muxrs2_outmux_2 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_766_ (
  .in1({ S193, S189 }),
  .out1({ S194 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_767_ (
  .in1({ new_datapath_muxrs2_outmux_2, new_datapath_muxrs2_outmux_1 }),
  .out1({ S195 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_768_ (
  .in1({ S195, S185 }),
  .out1({ S196 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_769_ (
  .in1({ S194, S184 }),
  .out1({ S197 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_770_ (
  .in1({ S196, new_controller_outflag_6 }),
  .out1({ S198 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_771_ (
  .in1({ S198 }),
  .out1({ S199 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_772_ (
  .in1({ S196, S3303 }),
  .out1({ S200 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_773_ (
  .in1({ S200 }),
  .out1({ S201 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_774_ (
  .in1({ S200, S199 }),
  .out1({ S202 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_775_ (
  .in1({ S201, S198 }),
  .out1({ S203 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_776_ (
  .in1({ S196, new_controller_407_B_2 }),
  .out1({ S204 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_777_ (
  .in1({ S204 }),
  .out1({ S205 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_778_ (
  .in1({ S196, S3292 }),
  .out1({ S206 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_779_ (
  .in1({ S206 }),
  .out1({ S207 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_780_ (
  .in1({ S206, S205 }),
  .out1({ S208 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_781_ (
  .in1({ S207, S204 }),
  .out1({ S209 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_782_ (
  .in1({ new_datapath_multdivunit_1697_B_14, new_datapath_multdivunit_1697_B_15 }),
  .out1({ S210 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_783_ (
  .in1({ S210 }),
  .out1({ S211 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_784_ (
  .in1({ S211, new_datapath_multdivunit_1697_B_13 }),
  .out1({ S212 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_785_ (
  .in1({ S212 }),
  .out1({ S213 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_786_ (
  .in1({ S213, new_datapath_multdivunit_1697_B_12 }),
  .out1({ S214 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_787_ (
  .in1({ S214 }),
  .out1({ S215 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_788_ (
  .in1({ S215, new_datapath_multdivunit_1697_B_11 }),
  .out1({ S216 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_789_ (
  .in1({ S214, S3445 }),
  .out1({ S217 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_790_ (
  .in1({ S217, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S218 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_791_ (
  .in1({ S218 }),
  .out1({ S219 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_792_ (
  .in1({ S219, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S220 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_793_ (
  .in1({ S220 }),
  .out1({ S221 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_794_ (
  .in1({ S221, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S222 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_795_ (
  .in1({ S222 }),
  .out1({ S223 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_796_ (
  .in1({ S197, S2614 }),
  .out1({ S224 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_797_ (
  .in1({ S196, new_controller_outflag_7 }),
  .out1({ S225 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_798_ (
  .in1({ S196, S3314 }),
  .out1({ S226 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_799_ (
  .in1({ S197, new_datapath_p2trf_7 }),
  .out1({ S227 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_800_ (
  .in1({ S226, S224 }),
  .out1({ S228 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_801_ (
  .in1({ S227, S225 }),
  .out1({ S229 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_802_ (
  .in1({ S229, S223 }),
  .out1({ S230 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_803_ (
  .in1({ S228, S222 }),
  .out1({ S231 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_804_ (
  .in1({ S231, S203 }),
  .out1({ S232 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_805_ (
  .in1({ S230, S202 }),
  .out1({ S233 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_806_ (
  .in1({ S233, S209 }),
  .out1({ S234 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_807_ (
  .in1({ S232, S208 }),
  .out1({ S235 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_808_ (
  .in1({ S196, new_controller_407_B_0 }),
  .out1({ S236 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_809_ (
  .in1({ S236 }),
  .out1({ S237 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_810_ (
  .in1({ S196, S3281 }),
  .out1({ S238 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_811_ (
  .in1({ S238 }),
  .out1({ S239 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_812_ (
  .in1({ S238, S237 }),
  .out1({ S240 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_813_ (
  .in1({ S239, S236 }),
  .out1({ S241 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_814_ (
  .in1({ S241, S235 }),
  .out1({ S242 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_815_ (
  .in1({ S240, S234 }),
  .out1({ S243 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_816_ (
  .in1({ S196, new_controller_outflag_3 }),
  .out1({ S244 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_817_ (
  .in1({ S244 }),
  .out1({ S245 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_818_ (
  .in1({ S196, S3270 }),
  .out1({ S246 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_819_ (
  .in1({ S246 }),
  .out1({ S247 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_820_ (
  .in1({ S246, S245 }),
  .out1({ S248 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_821_ (
  .in1({ S247, S244 }),
  .out1({ S249 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_822_ (
  .in1({ S249, S243 }),
  .out1({ S250 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_823_ (
  .in1({ S248, S242 }),
  .out1({ S251 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_824_ (
  .in1({ S196, new_controller_outflag_2 }),
  .out1({ S252 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_825_ (
  .in1({ S252 }),
  .out1({ S253 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_826_ (
  .in1({ S196, S3259 }),
  .out1({ S254 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_827_ (
  .in1({ S254 }),
  .out1({ S255 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_828_ (
  .in1({ S254, S253 }),
  .out1({ S256 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_829_ (
  .in1({ S255, S252 }),
  .out1({ S257 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_830_ (
  .in1({ S257, S251 }),
  .out1({ S258 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_831_ (
  .in1({ S256, S250 }),
  .out1({ S259 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_832_ (
  .in1({ S196, new_controller_outflag_1 }),
  .out1({ S260 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_833_ (
  .in1({ S260 }),
  .out1({ S261 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_834_ (
  .in1({ S196, S3248 }),
  .out1({ S262 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_835_ (
  .in1({ S262 }),
  .out1({ S263 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_836_ (
  .in1({ S262, S261 }),
  .out1({ S264 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_837_ (
  .in1({ S263, S260 }),
  .out1({ S265 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_838_ (
  .in1({ S196, new_controller_outflag_0 }),
  .out1({ S266 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_839_ (
  .in1({ S266 }),
  .out1({ S267 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_840_ (
  .in1({ S196, S3237 }),
  .out1({ S268 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_841_ (
  .in1({ S268 }),
  .out1({ S269 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_842_ (
  .in1({ S268, S267 }),
  .out1({ S270 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_843_ (
  .in1({ S269, S266 }),
  .out1({ S271 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_844_ (
  .in1({ S265, S259 }),
  .out1({ S272 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_845_ (
  .in1({ S264, S258 }),
  .out1({ S273 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_846_ (
  .in1({ S273, S270 }),
  .out1({ S274 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_847_ (
  .in1({ S272, S271 }),
  .out1({ S275 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_848_ (
  .in1({ S274, S3401 }),
  .out1({ S276 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_849_ (
  .in1({ S275, new_datapath_addsubunit_in1_15 }),
  .out1({ S277 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_850_ (
  .in1({ S277, S265 }),
  .out1({ S278 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_851_ (
  .in1({ S276, S264 }),
  .out1({ S279 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_852_ (
  .in1({ S264, new_datapath_addsubunit_in1_15 }),
  .out1({ S280 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_853_ (
  .in1({ S265, S3401 }),
  .out1({ S281 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_854_ (
  .in1({ S280, S278 }),
  .out1({ S282 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_855_ (
  .in1({ S281, S279 }),
  .out1({ S283 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_856_ (
  .in1({ S270, new_datapath_addsubunit_in1_14 }),
  .out1({ S284 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_857_ (
  .in1({ S271, S3390 }),
  .out1({ S285 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_858_ (
  .in1({ S284, S283 }),
  .out1({ S286 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_859_ (
  .in1({ S285, S282 }),
  .out1({ S287 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_860_ (
  .in1({ S286, S278 }),
  .out1({ S288 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_861_ (
  .in1({ S287, S279 }),
  .out1({ S289 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_862_ (
  .in1({ S288, S259 }),
  .out1({ S290 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_863_ (
  .in1({ S289, S258 }),
  .out1({ S291 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_864_ (
  .in1({ S285, S282 }),
  .out1({ S292 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_865_ (
  .in1({ S292, S286 }),
  .out1({ S293 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_866_ (
  .in1({ S290, S277 }),
  .out1({ S294 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_867_ (
  .in1({ S291, S276 }),
  .out1({ S295 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_868_ (
  .in1({ S293, S290 }),
  .out1({ S296 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_869_ (
  .in1({ S296 }),
  .out1({ S297 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_870_ (
  .in1({ S296, S295 }),
  .out1({ S298 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_871_ (
  .in1({ S297, S294 }),
  .out1({ S299 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_872_ (
  .in1({ S291, S270 }),
  .out1({ S300 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_873_ (
  .in1({ S290, S271 }),
  .out1({ S301 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_874_ (
  .in1({ S300, S3390 }),
  .out1({ S302 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_875_ (
  .in1({ S301, new_datapath_addsubunit_in1_14 }),
  .out1({ S303 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_876_ (
  .in1({ S303, S265 }),
  .out1({ S304 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_877_ (
  .in1({ S302, S264 }),
  .out1({ S305 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_878_ (
  .in1({ S302, S264 }),
  .out1({ S306 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_879_ (
  .in1({ S303, S265 }),
  .out1({ S307 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_880_ (
  .in1({ S306, S304 }),
  .out1({ S308 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_881_ (
  .in1({ S307, S305 }),
  .out1({ S309 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_882_ (
  .in1({ S270, new_datapath_addsubunit_in1_13 }),
  .out1({ S310 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_883_ (
  .in1({ S271, S3379 }),
  .out1({ S311 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_884_ (
  .in1({ S310, S309 }),
  .out1({ S312 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_885_ (
  .in1({ S311, S308 }),
  .out1({ S313 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_886_ (
  .in1({ S312, S304 }),
  .out1({ S314 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_887_ (
  .in1({ S313, S305 }),
  .out1({ S315 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_888_ (
  .in1({ S257, S250 }),
  .out1({ S316 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_889_ (
  .in1({ S316, S314 }),
  .out1({ S317 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_890_ (
  .in1({ S314, S258 }),
  .out1({ S318 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_891_ (
  .in1({ S318, S298 }),
  .out1({ S319 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_892_ (
  .in1({ S317, S299 }),
  .out1({ S320 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_893_ (
  .in1({ S319, S317 }),
  .out1({ S321 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_894_ (
  .in1({ S320, S318 }),
  .out1({ S322 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_895_ (
  .in1({ S299, S257 }),
  .out1({ S323 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_896_ (
  .in1({ S298, S256 }),
  .out1({ S324 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_897_ (
  .in1({ S323, S315 }),
  .out1({ S325 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_898_ (
  .in1({ S324, S314 }),
  .out1({ S326 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_899_ (
  .in1({ S256, new_datapath_addsubunit_in1_15 }),
  .out1({ S327 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_900_ (
  .in1({ S257, S3401 }),
  .out1({ S328 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_901_ (
  .in1({ S327, S251 }),
  .out1({ S329 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_902_ (
  .in1({ S328, S250 }),
  .out1({ S330 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_903_ (
  .in1({ S330, S325 }),
  .out1({ S331 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_904_ (
  .in1({ S329, S326 }),
  .out1({ S332 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_905_ (
  .in1({ S310, S309 }),
  .out1({ S333 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_906_ (
  .in1({ S333, S313 }),
  .out1({ S334 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_907_ (
  .in1({ S331, S303 }),
  .out1({ S335 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_908_ (
  .in1({ S332, S302 }),
  .out1({ S336 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_909_ (
  .in1({ S334, S332 }),
  .out1({ S337 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_910_ (
  .in1({ S337 }),
  .out1({ S338 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_911_ (
  .in1({ S338, S336 }),
  .out1({ S339 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_912_ (
  .in1({ S337, S335 }),
  .out1({ S340 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_913_ (
  .in1({ S340, S257 }),
  .out1({ S341 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_914_ (
  .in1({ S339, S256 }),
  .out1({ S342 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_915_ (
  .in1({ S339, S256 }),
  .out1({ S343 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_916_ (
  .in1({ S340, S257 }),
  .out1({ S344 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_917_ (
  .in1({ S343, S341 }),
  .out1({ S345 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_918_ (
  .in1({ S344, S342 }),
  .out1({ S346 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_919_ (
  .in1({ S331, new_datapath_addsubunit_in1_13 }),
  .out1({ S347 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_920_ (
  .in1({ S332, S3379 }),
  .out1({ S348 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_921_ (
  .in1({ S271, new_datapath_addsubunit_in1_13 }),
  .out1({ S349 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_922_ (
  .in1({ S349 }),
  .out1({ S350 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_923_ (
  .in1({ S270, S3379 }),
  .out1({ S351 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_924_ (
  .in1({ S271, new_datapath_addsubunit_in1_13 }),
  .out1({ S352 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_925_ (
  .in1({ S352, S350 }),
  .out1({ S353 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_926_ (
  .in1({ S351, S349 }),
  .out1({ S354 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_927_ (
  .in1({ S354, S332 }),
  .out1({ S355 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_928_ (
  .in1({ S353, S331 }),
  .out1({ S356 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_929_ (
  .in1({ S355, S347 }),
  .out1({ S357 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_930_ (
  .in1({ S356, S348 }),
  .out1({ S358 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_931_ (
  .in1({ S358, S265 }),
  .out1({ S359 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_932_ (
  .in1({ S357, S264 }),
  .out1({ S360 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_933_ (
  .in1({ S270, new_datapath_addsubunit_in1_12 }),
  .out1({ S361 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_934_ (
  .in1({ S271, S3368 }),
  .out1({ S362 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_935_ (
  .in1({ S357, S264 }),
  .out1({ S363 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_936_ (
  .in1({ S358, S265 }),
  .out1({ S364 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_937_ (
  .in1({ S363, S359 }),
  .out1({ S365 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_938_ (
  .in1({ S364, S360 }),
  .out1({ S366 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_939_ (
  .in1({ S366, S361 }),
  .out1({ S367 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_940_ (
  .in1({ S365, S362 }),
  .out1({ S368 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_941_ (
  .in1({ S367, S359 }),
  .out1({ S369 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_942_ (
  .in1({ S368, S360 }),
  .out1({ S370 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_943_ (
  .in1({ S369, S346 }),
  .out1({ S371 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_944_ (
  .in1({ S370, S345 }),
  .out1({ S372 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_945_ (
  .in1({ S371, S341 }),
  .out1({ S373 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_946_ (
  .in1({ S372, S342 }),
  .out1({ S374 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_947_ (
  .in1({ S373, S249 }),
  .out1({ S375 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_948_ (
  .in1({ S374, S248 }),
  .out1({ S376 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_949_ (
  .in1({ S374, S248 }),
  .out1({ S377 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_950_ (
  .in1({ S373, S249 }),
  .out1({ S378 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_951_ (
  .in1({ S377, S243 }),
  .out1({ S379 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_952_ (
  .in1({ S378, S242 }),
  .out1({ S380 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_953_ (
  .in1({ S380, S375 }),
  .out1({ S381 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_954_ (
  .in1({ S381, S322 }),
  .out1({ S382 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_955_ (
  .in1({ S382 }),
  .out1({ S383 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_956_ (
  .in1({ S383, S241 }),
  .out1({ S384 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_957_ (
  .in1({ S382, S240 }),
  .out1({ S385 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_958_ (
  .in1({ S321, S240 }),
  .out1({ S386 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_959_ (
  .in1({ S322, S241 }),
  .out1({ S387 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_960_ (
  .in1({ S386, S384 }),
  .out1({ S388 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_961_ (
  .in1({ S387, S385 }),
  .out1({ S389 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_962_ (
  .in1({ S375, S321 }),
  .out1({ S390 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_963_ (
  .in1({ S376, S322 }),
  .out1({ S391 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_964_ (
  .in1({ S390, S380 }),
  .out1({ S392 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_965_ (
  .in1({ S391, S379 }),
  .out1({ S393 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_966_ (
  .in1({ S370, S345 }),
  .out1({ S394 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_967_ (
  .in1({ S369, S346 }),
  .out1({ S395 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_968_ (
  .in1({ S394, S371 }),
  .out1({ S396 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_969_ (
  .in1({ S395, S372 }),
  .out1({ S397 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_970_ (
  .in1({ S396, S393 }),
  .out1({ S398 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_971_ (
  .in1({ S397, S392 }),
  .out1({ S399 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_972_ (
  .in1({ S392, S339 }),
  .out1({ S400 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_973_ (
  .in1({ S393, S340 }),
  .out1({ S401 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_974_ (
  .in1({ S400, S398 }),
  .out1({ S402 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_975_ (
  .in1({ S401, S399 }),
  .out1({ S403 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_976_ (
  .in1({ S403, S249 }),
  .out1({ S404 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_977_ (
  .in1({ S402, S248 }),
  .out1({ S405 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_978_ (
  .in1({ S402, S248 }),
  .out1({ S406 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_979_ (
  .in1({ S403, S249 }),
  .out1({ S407 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_980_ (
  .in1({ S406, S404 }),
  .out1({ S408 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_981_ (
  .in1({ S407, S405 }),
  .out1({ S409 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_982_ (
  .in1({ S365, S362 }),
  .out1({ S410 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_983_ (
  .in1({ S366, S361 }),
  .out1({ S411 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_984_ (
  .in1({ S410, S367 }),
  .out1({ S412 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_985_ (
  .in1({ S411, S368 }),
  .out1({ S413 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_986_ (
  .in1({ S413, S393 }),
  .out1({ S414 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_987_ (
  .in1({ S412, S392 }),
  .out1({ S415 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_988_ (
  .in1({ S392, S358 }),
  .out1({ S416 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_989_ (
  .in1({ S393, S357 }),
  .out1({ S417 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_990_ (
  .in1({ S416, S414 }),
  .out1({ S418 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_991_ (
  .in1({ S417, S415 }),
  .out1({ S419 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_992_ (
  .in1({ S418, S257 }),
  .out1({ S420 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_993_ (
  .in1({ S419, S256 }),
  .out1({ S421 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_994_ (
  .in1({ S419, S256 }),
  .out1({ S422 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_995_ (
  .in1({ S418, S257 }),
  .out1({ S423 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_996_ (
  .in1({ S422, S420 }),
  .out1({ S424 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_997_ (
  .in1({ S423, S421 }),
  .out1({ S425 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_998_ (
  .in1({ S271, S3368 }),
  .out1({ S426 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_999_ (
  .in1({ S270, new_datapath_addsubunit_in1_12 }),
  .out1({ S427 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1000_ (
  .in1({ S426, S361 }),
  .out1({ S428 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1001_ (
  .in1({ S427, S362 }),
  .out1({ S429 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1002_ (
  .in1({ S428, S393 }),
  .out1({ S430 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1003_ (
  .in1({ S429, S392 }),
  .out1({ S431 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1004_ (
  .in1({ S392, S3368 }),
  .out1({ S432 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1005_ (
  .in1({ S393, new_datapath_addsubunit_in1_12 }),
  .out1({ S433 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1006_ (
  .in1({ S432, S430 }),
  .out1({ S434 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1007_ (
  .in1({ S433, S431 }),
  .out1({ S435 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1008_ (
  .in1({ S434, S265 }),
  .out1({ S436 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1009_ (
  .in1({ S435, S264 }),
  .out1({ S437 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1010_ (
  .in1({ S435, S264 }),
  .out1({ S438 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1011_ (
  .in1({ S434, S265 }),
  .out1({ S439 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1012_ (
  .in1({ S438, S436 }),
  .out1({ S440 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1013_ (
  .in1({ S439, S437 }),
  .out1({ S441 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1014_ (
  .in1({ S270, new_datapath_addsubunit_in1_11 }),
  .out1({ S442 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1015_ (
  .in1({ S271, S3357 }),
  .out1({ S443 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1016_ (
  .in1({ S442, S441 }),
  .out1({ S444 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1017_ (
  .in1({ S443, S440 }),
  .out1({ S445 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1018_ (
  .in1({ S444, S436 }),
  .out1({ S446 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1019_ (
  .in1({ S445, S437 }),
  .out1({ S447 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1020_ (
  .in1({ S446, S425 }),
  .out1({ S448 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1021_ (
  .in1({ S447, S424 }),
  .out1({ S449 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1022_ (
  .in1({ S448, S420 }),
  .out1({ S450 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1023_ (
  .in1({ S449, S421 }),
  .out1({ S451 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1024_ (
  .in1({ S450, S409 }),
  .out1({ S452 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1025_ (
  .in1({ S451, S408 }),
  .out1({ S453 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1026_ (
  .in1({ S452, S404 }),
  .out1({ S454 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1027_ (
  .in1({ S453, S405 }),
  .out1({ S455 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1028_ (
  .in1({ S454, S389 }),
  .out1({ S456 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1029_ (
  .in1({ S455, S388 }),
  .out1({ S457 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1030_ (
  .in1({ S456, S384 }),
  .out1({ S458 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1031_ (
  .in1({ S457, S385 }),
  .out1({ S459 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1032_ (
  .in1({ S458, S235 }),
  .out1({ S460 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1033_ (
  .in1({ S459, S234 }),
  .out1({ S461 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1034_ (
  .in1({ S461, S382 }),
  .out1({ S462 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1035_ (
  .in1({ S462, S296 }),
  .out1({ S463 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1036_ (
  .in1({ S463 }),
  .out1({ S464 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1037_ (
  .in1({ S451, S408 }),
  .out1({ S465 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1038_ (
  .in1({ S465, S452 }),
  .out1({ S466 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1039_ (
  .in1({ S466, S461 }),
  .out1({ S467 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1040_ (
  .in1({ S467 }),
  .out1({ S468 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1041_ (
  .in1({ S460, S402 }),
  .out1({ S469 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1042_ (
  .in1({ S461, S403 }),
  .out1({ S470 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1043_ (
  .in1({ S469, S467 }),
  .out1({ S471 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1044_ (
  .in1({ S470, S468 }),
  .out1({ S472 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1045_ (
  .in1({ S472, S241 }),
  .out1({ S473 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1046_ (
  .in1({ S471, S240 }),
  .out1({ S474 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1047_ (
  .in1({ S471, S240 }),
  .out1({ S475 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1048_ (
  .in1({ S472, S241 }),
  .out1({ S476 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1049_ (
  .in1({ S475, S473 }),
  .out1({ S477 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1050_ (
  .in1({ S476, S474 }),
  .out1({ S478 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1051_ (
  .in1({ S447, S424 }),
  .out1({ S479 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1052_ (
  .in1({ S479, S448 }),
  .out1({ S480 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1053_ (
  .in1({ S480, S461 }),
  .out1({ S481 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1054_ (
  .in1({ S481 }),
  .out1({ S482 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1055_ (
  .in1({ S460, S419 }),
  .out1({ S483 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1056_ (
  .in1({ S461, S418 }),
  .out1({ S484 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1057_ (
  .in1({ S483, S481 }),
  .out1({ S485 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1058_ (
  .in1({ S484, S482 }),
  .out1({ S486 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1059_ (
  .in1({ S486, S249 }),
  .out1({ S487 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1060_ (
  .in1({ S485, S248 }),
  .out1({ S488 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1061_ (
  .in1({ S485, S248 }),
  .out1({ S489 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1062_ (
  .in1({ S486, S249 }),
  .out1({ S490 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1063_ (
  .in1({ S489, S487 }),
  .out1({ S491 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1064_ (
  .in1({ S490, S488 }),
  .out1({ S492 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1065_ (
  .in1({ S442, S441 }),
  .out1({ S493 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1066_ (
  .in1({ S493, S445 }),
  .out1({ S494 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1067_ (
  .in1({ S494, S461 }),
  .out1({ S495 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1068_ (
  .in1({ S495 }),
  .out1({ S496 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1069_ (
  .in1({ S461, S435 }),
  .out1({ S497 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1070_ (
  .in1({ S497 }),
  .out1({ S498 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1071_ (
  .in1({ S498, S495 }),
  .out1({ S499 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1072_ (
  .in1({ S497, S496 }),
  .out1({ S500 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1073_ (
  .in1({ S499, S257 }),
  .out1({ S501 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1074_ (
  .in1({ S500, S256 }),
  .out1({ S502 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1075_ (
  .in1({ S500, S256 }),
  .out1({ S503 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1076_ (
  .in1({ S499, S257 }),
  .out1({ S504 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1077_ (
  .in1({ S503, S501 }),
  .out1({ S505 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1078_ (
  .in1({ S504, S502 }),
  .out1({ S506 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1079_ (
  .in1({ S460, new_datapath_addsubunit_in1_11 }),
  .out1({ S507 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1080_ (
  .in1({ S461, S3357 }),
  .out1({ S508 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1081_ (
  .in1({ S271, new_datapath_addsubunit_in1_11 }),
  .out1({ S509 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1082_ (
  .in1({ S509 }),
  .out1({ S510 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1083_ (
  .in1({ S270, S3357 }),
  .out1({ S511 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1084_ (
  .in1({ S271, new_datapath_addsubunit_in1_11 }),
  .out1({ S512 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1085_ (
  .in1({ S512, S510 }),
  .out1({ S513 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1086_ (
  .in1({ S511, S509 }),
  .out1({ S514 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1087_ (
  .in1({ S514, S461 }),
  .out1({ S515 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1088_ (
  .in1({ S513, S460 }),
  .out1({ S516 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1089_ (
  .in1({ S515, S507 }),
  .out1({ S517 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1090_ (
  .in1({ S516, S508 }),
  .out1({ S518 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1091_ (
  .in1({ S518, S265 }),
  .out1({ S519 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1092_ (
  .in1({ S517, S264 }),
  .out1({ S520 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1093_ (
  .in1({ S270, new_datapath_addsubunit_in1_10 }),
  .out1({ S521 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1094_ (
  .in1({ S271, S3346 }),
  .out1({ S522 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1095_ (
  .in1({ S517, S264 }),
  .out1({ S523 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1096_ (
  .in1({ S518, S265 }),
  .out1({ S524 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1097_ (
  .in1({ S523, S519 }),
  .out1({ S525 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1098_ (
  .in1({ S524, S520 }),
  .out1({ S526 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1099_ (
  .in1({ S526, S521 }),
  .out1({ S527 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1100_ (
  .in1({ S525, S522 }),
  .out1({ S528 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1101_ (
  .in1({ S527, S519 }),
  .out1({ S529 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1102_ (
  .in1({ S528, S520 }),
  .out1({ S530 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1103_ (
  .in1({ S529, S506 }),
  .out1({ S531 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1104_ (
  .in1({ S530, S505 }),
  .out1({ S532 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1105_ (
  .in1({ S531, S501 }),
  .out1({ S533 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1106_ (
  .in1({ S532, S502 }),
  .out1({ S534 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1107_ (
  .in1({ S533, S492 }),
  .out1({ S535 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1108_ (
  .in1({ S534, S491 }),
  .out1({ S536 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1109_ (
  .in1({ S535, S487 }),
  .out1({ S537 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1110_ (
  .in1({ S536, S488 }),
  .out1({ S538 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1111_ (
  .in1({ S537, S478 }),
  .out1({ S539 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1112_ (
  .in1({ S538, S477 }),
  .out1({ S540 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1113_ (
  .in1({ S539, S473 }),
  .out1({ S541 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1114_ (
  .in1({ S540, S474 }),
  .out1({ S542 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1115_ (
  .in1({ S232, S209 }),
  .out1({ S543 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1116_ (
  .in1({ S543, S542 }),
  .out1({ S544 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1117_ (
  .in1({ S541, S235 }),
  .out1({ S545 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1118_ (
  .in1({ S545, S544 }),
  .out1({ S546 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1119_ (
  .in1({ S546, S463 }),
  .out1({ S547 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1120_ (
  .in1({ S464, S209 }),
  .out1({ S548 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1121_ (
  .in1({ S463, S208 }),
  .out1({ S549 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1122_ (
  .in1({ S548, S542 }),
  .out1({ S550 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1123_ (
  .in1({ S549, S541 }),
  .out1({ S551 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1124_ (
  .in1({ S463, S208 }),
  .out1({ S552 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1125_ (
  .in1({ S464, S209 }),
  .out1({ S553 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1126_ (
  .in1({ S552, S233 }),
  .out1({ S554 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1127_ (
  .in1({ S553, S232 }),
  .out1({ S555 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1128_ (
  .in1({ S555, S550 }),
  .out1({ S556 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1129_ (
  .in1({ S554, S551 }),
  .out1({ S557 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1130_ (
  .in1({ S537, S478 }),
  .out1({ S558 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1131_ (
  .in1({ S558, S540 }),
  .out1({ S559 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1132_ (
  .in1({ S559, S556 }),
  .out1({ S560 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1133_ (
  .in1({ S557, S472 }),
  .out1({ S561 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1134_ (
  .in1({ S561, S560 }),
  .out1({ S562 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1135_ (
  .in1({ S562 }),
  .out1({ S563 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1136_ (
  .in1({ S562, S209 }),
  .out1({ S564 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1137_ (
  .in1({ S563, S208 }),
  .out1({ S565 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1138_ (
  .in1({ S563, S208 }),
  .out1({ S566 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1139_ (
  .in1({ S566, S564 }),
  .out1({ S567 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1140_ (
  .in1({ S567 }),
  .out1({ S568 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1141_ (
  .in1({ S533, S492 }),
  .out1({ S569 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1142_ (
  .in1({ S569, S536 }),
  .out1({ S570 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1143_ (
  .in1({ S570, S556 }),
  .out1({ S571 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1144_ (
  .in1({ S571 }),
  .out1({ S572 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1145_ (
  .in1({ S556, S485 }),
  .out1({ S573 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1146_ (
  .in1({ S573 }),
  .out1({ S574 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1147_ (
  .in1({ S573, S572 }),
  .out1({ S575 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1148_ (
  .in1({ S574, S571 }),
  .out1({ S576 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1149_ (
  .in1({ S576, S241 }),
  .out1({ S577 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1150_ (
  .in1({ S575, S240 }),
  .out1({ S578 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1151_ (
  .in1({ S575, S240 }),
  .out1({ S579 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1152_ (
  .in1({ S576, S241 }),
  .out1({ S580 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1153_ (
  .in1({ S579, S577 }),
  .out1({ S581 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1154_ (
  .in1({ S580, S578 }),
  .out1({ S582 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1155_ (
  .in1({ S529, S506 }),
  .out1({ S583 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1156_ (
  .in1({ S583, S532 }),
  .out1({ S584 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1157_ (
  .in1({ S584, S556 }),
  .out1({ S585 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1158_ (
  .in1({ S557, S499 }),
  .out1({ S586 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1159_ (
  .in1({ S586, S585 }),
  .out1({ S587 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1160_ (
  .in1({ S587 }),
  .out1({ S588 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1161_ (
  .in1({ S587, S249 }),
  .out1({ S589 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1162_ (
  .in1({ S588, S248 }),
  .out1({ S590 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1163_ (
  .in1({ S587, S249 }),
  .out1({ S591 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1164_ (
  .in1({ S591 }),
  .out1({ S592 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1165_ (
  .in1({ S592, S589 }),
  .out1({ S593 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1166_ (
  .in1({ S593 }),
  .out1({ S594 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1167_ (
  .in1({ S525, S522 }),
  .out1({ S595 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1168_ (
  .in1({ S526, S521 }),
  .out1({ S596 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1169_ (
  .in1({ S595, S527 }),
  .out1({ S597 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1170_ (
  .in1({ S596, S528 }),
  .out1({ S598 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1171_ (
  .in1({ S598, S557 }),
  .out1({ S599 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1172_ (
  .in1({ S597, S556 }),
  .out1({ S600 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1173_ (
  .in1({ S556, S518 }),
  .out1({ S601 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1174_ (
  .in1({ S557, S517 }),
  .out1({ S602 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1175_ (
  .in1({ S601, S599 }),
  .out1({ S603 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1176_ (
  .in1({ S602, S600 }),
  .out1({ S604 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1177_ (
  .in1({ S603, S257 }),
  .out1({ S605 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1178_ (
  .in1({ S604, S256 }),
  .out1({ S606 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1179_ (
  .in1({ S604, S256 }),
  .out1({ S607 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1180_ (
  .in1({ S603, S257 }),
  .out1({ S608 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1181_ (
  .in1({ S607, S605 }),
  .out1({ S609 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1182_ (
  .in1({ S608, S606 }),
  .out1({ S610 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1183_ (
  .in1({ S556, new_datapath_addsubunit_in1_10 }),
  .out1({ S611 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1184_ (
  .in1({ S557, S3346 }),
  .out1({ S612 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1185_ (
  .in1({ S271, S3346 }),
  .out1({ S613 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1186_ (
  .in1({ S270, new_datapath_addsubunit_in1_10 }),
  .out1({ S614 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1187_ (
  .in1({ S613, S521 }),
  .out1({ S615 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1188_ (
  .in1({ S614, S522 }),
  .out1({ S616 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1189_ (
  .in1({ S616, S557 }),
  .out1({ S617 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1190_ (
  .in1({ S615, S556 }),
  .out1({ S618 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1191_ (
  .in1({ S617, S611 }),
  .out1({ S619 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1192_ (
  .in1({ S618, S612 }),
  .out1({ S620 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1193_ (
  .in1({ S620, S265 }),
  .out1({ S621 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1194_ (
  .in1({ S619, S264 }),
  .out1({ S622 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1195_ (
  .in1({ S619, S264 }),
  .out1({ S623 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1196_ (
  .in1({ S620, S265 }),
  .out1({ S624 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1197_ (
  .in1({ S623, S621 }),
  .out1({ S625 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1198_ (
  .in1({ S624, S622 }),
  .out1({ S626 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1199_ (
  .in1({ S270, new_datapath_addsubunit_in1_9 }),
  .out1({ S627 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1200_ (
  .in1({ S271, S3336 }),
  .out1({ S628 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1201_ (
  .in1({ S627, S626 }),
  .out1({ S629 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1202_ (
  .in1({ S628, S625 }),
  .out1({ S630 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1203_ (
  .in1({ S629, S621 }),
  .out1({ S631 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1204_ (
  .in1({ S630, S622 }),
  .out1({ S632 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1205_ (
  .in1({ S631, S610 }),
  .out1({ S633 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1206_ (
  .in1({ S632, S609 }),
  .out1({ S634 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1207_ (
  .in1({ S633, S605 }),
  .out1({ S635 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1208_ (
  .in1({ S634, S606 }),
  .out1({ S636 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1209_ (
  .in1({ S635, S594 }),
  .out1({ S637 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1210_ (
  .in1({ S636, S593 }),
  .out1({ S638 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1211_ (
  .in1({ S637, S589 }),
  .out1({ S639 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1212_ (
  .in1({ S638, S590 }),
  .out1({ S640 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1213_ (
  .in1({ S639, S582 }),
  .out1({ S641 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1214_ (
  .in1({ S640, S581 }),
  .out1({ S642 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1215_ (
  .in1({ S641, S577 }),
  .out1({ S643 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1216_ (
  .in1({ S642, S578 }),
  .out1({ S644 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1217_ (
  .in1({ S643, S568 }),
  .out1({ S645 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1218_ (
  .in1({ S644, S567 }),
  .out1({ S646 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1219_ (
  .in1({ S645, S564 }),
  .out1({ S647 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1220_ (
  .in1({ S646, S565 }),
  .out1({ S648 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1221_ (
  .in1({ S230, S203 }),
  .out1({ S649 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1222_ (
  .in1({ S647, S232 }),
  .out1({ S650 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1223_ (
  .in1({ S649, S647 }),
  .out1({ S651 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1224_ (
  .in1({ S651, S547 }),
  .out1({ S652 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1225_ (
  .in1({ S652, S650 }),
  .out1({ S653 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1226_ (
  .in1({ S653 }),
  .out1({ S654 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1227_ (
  .in1({ S547, S203 }),
  .out1({ S655 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1228_ (
  .in1({ S655 }),
  .out1({ S656 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1229_ (
  .in1({ S655, S648 }),
  .out1({ S657 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1230_ (
  .in1({ S656, S647 }),
  .out1({ S658 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1231_ (
  .in1({ S463, S202 }),
  .out1({ S659 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1232_ (
  .in1({ S464, S203 }),
  .out1({ S660 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1233_ (
  .in1({ S659, S231 }),
  .out1({ S661 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1234_ (
  .in1({ S660, S230 }),
  .out1({ S662 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1235_ (
  .in1({ S662, S657 }),
  .out1({ S663 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1236_ (
  .in1({ S661, S658 }),
  .out1({ S664 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1237_ (
  .in1({ S644, S567 }),
  .out1({ S665 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1238_ (
  .in1({ S665, S645 }),
  .out1({ S666 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1239_ (
  .in1({ S666, S664 }),
  .out1({ S667 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1240_ (
  .in1({ S667 }),
  .out1({ S668 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1241_ (
  .in1({ S664, S562 }),
  .out1({ S669 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1242_ (
  .in1({ S669 }),
  .out1({ S670 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1243_ (
  .in1({ S670, S667 }),
  .out1({ S671 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1244_ (
  .in1({ S669, S668 }),
  .out1({ S672 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1245_ (
  .in1({ S672, S203 }),
  .out1({ S673 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1246_ (
  .in1({ S671, S202 }),
  .out1({ S674 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1247_ (
  .in1({ S671, S202 }),
  .out1({ S675 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1248_ (
  .in1({ S672, S203 }),
  .out1({ S676 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1249_ (
  .in1({ S675, S673 }),
  .out1({ S677 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1250_ (
  .in1({ S676, S674 }),
  .out1({ S678 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1251_ (
  .in1({ S639, S582 }),
  .out1({ S679 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1252_ (
  .in1({ S679 }),
  .out1({ S680 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1253_ (
  .in1({ S680, S641 }),
  .out1({ S681 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1254_ (
  .in1({ S681, S664 }),
  .out1({ S682 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1255_ (
  .in1({ S682 }),
  .out1({ S683 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1256_ (
  .in1({ S663, S575 }),
  .out1({ S684 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1257_ (
  .in1({ S664, S576 }),
  .out1({ S685 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1258_ (
  .in1({ S684, S682 }),
  .out1({ S686 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1259_ (
  .in1({ S685, S683 }),
  .out1({ S687 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1260_ (
  .in1({ S687, S209 }),
  .out1({ S688 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1261_ (
  .in1({ S686, S208 }),
  .out1({ S689 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1262_ (
  .in1({ S686, S208 }),
  .out1({ S690 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1263_ (
  .in1({ S687, S209 }),
  .out1({ S691 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1264_ (
  .in1({ S690, S688 }),
  .out1({ S692 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1265_ (
  .in1({ S691, S689 }),
  .out1({ S693 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1266_ (
  .in1({ S635, S594 }),
  .out1({ S694 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1267_ (
  .in1({ S694, S638 }),
  .out1({ S695 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1268_ (
  .in1({ S695, S663 }),
  .out1({ S696 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1269_ (
  .in1({ S664, S587 }),
  .out1({ S697 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1270_ (
  .in1({ S697, S696 }),
  .out1({ S698 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1271_ (
  .in1({ S698 }),
  .out1({ S699 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1272_ (
  .in1({ S698, S241 }),
  .out1({ S700 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1273_ (
  .in1({ S699, S240 }),
  .out1({ S701 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1274_ (
  .in1({ S698, S241 }),
  .out1({ S702 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1275_ (
  .in1({ S702 }),
  .out1({ S703 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1276_ (
  .in1({ S703, S700 }),
  .out1({ S704 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1277_ (
  .in1({ S704 }),
  .out1({ S705 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1278_ (
  .in1({ S631, S610 }),
  .out1({ S706 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1279_ (
  .in1({ S706, S634 }),
  .out1({ S707 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1280_ (
  .in1({ S707, S663 }),
  .out1({ S708 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1281_ (
  .in1({ S664, S603 }),
  .out1({ S709 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1282_ (
  .in1({ S709, S708 }),
  .out1({ S710 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1283_ (
  .in1({ S710 }),
  .out1({ S711 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1284_ (
  .in1({ S710, S249 }),
  .out1({ S712 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1285_ (
  .in1({ S711, S248 }),
  .out1({ S713 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1286_ (
  .in1({ S710, S249 }),
  .out1({ S714 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1287_ (
  .in1({ S714 }),
  .out1({ S715 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1288_ (
  .in1({ S715, S712 }),
  .out1({ S716 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1289_ (
  .in1({ S716 }),
  .out1({ S717 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1290_ (
  .in1({ S628, S625 }),
  .out1({ S718 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1291_ (
  .in1({ S718, S629 }),
  .out1({ S719 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1292_ (
  .in1({ S719, S664 }),
  .out1({ S720 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1293_ (
  .in1({ S720 }),
  .out1({ S721 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1294_ (
  .in1({ S663, S619 }),
  .out1({ S722 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1295_ (
  .in1({ S664, S620 }),
  .out1({ S723 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1296_ (
  .in1({ S722, S720 }),
  .out1({ S724 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1297_ (
  .in1({ S723, S721 }),
  .out1({ S725 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1298_ (
  .in1({ S725, S257 }),
  .out1({ S726 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1299_ (
  .in1({ S724, S256 }),
  .out1({ S727 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1300_ (
  .in1({ S724, S256 }),
  .out1({ S728 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1301_ (
  .in1({ S725, S257 }),
  .out1({ S729 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1302_ (
  .in1({ S728, S726 }),
  .out1({ S730 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1303_ (
  .in1({ S729, S727 }),
  .out1({ S731 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1304_ (
  .in1({ S663, new_datapath_addsubunit_in1_9 }),
  .out1({ S732 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1305_ (
  .in1({ S664, S3336 }),
  .out1({ S733 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1306_ (
  .in1({ S271, new_datapath_addsubunit_in1_9 }),
  .out1({ S734 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1307_ (
  .in1({ S734 }),
  .out1({ S735 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1308_ (
  .in1({ S270, S3336 }),
  .out1({ S736 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1309_ (
  .in1({ S271, new_datapath_addsubunit_in1_9 }),
  .out1({ S737 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1310_ (
  .in1({ S737, S735 }),
  .out1({ S738 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1311_ (
  .in1({ S736, S734 }),
  .out1({ S739 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1312_ (
  .in1({ S739, S664 }),
  .out1({ S740 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1313_ (
  .in1({ S738, S663 }),
  .out1({ S741 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1314_ (
  .in1({ S740, S732 }),
  .out1({ S742 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1315_ (
  .in1({ S741, S733 }),
  .out1({ S743 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1316_ (
  .in1({ S743, S265 }),
  .out1({ S744 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1317_ (
  .in1({ S742, S264 }),
  .out1({ S745 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1318_ (
  .in1({ S270, new_datapath_addsubunit_in1_8 }),
  .out1({ S746 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1319_ (
  .in1({ S271, S3325 }),
  .out1({ S747 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1320_ (
  .in1({ S742, S264 }),
  .out1({ S748 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1321_ (
  .in1({ S743, S265 }),
  .out1({ S749 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1322_ (
  .in1({ S748, S744 }),
  .out1({ S750 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1323_ (
  .in1({ S749, S745 }),
  .out1({ S751 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1324_ (
  .in1({ S751, S746 }),
  .out1({ S752 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1325_ (
  .in1({ S750, S747 }),
  .out1({ S753 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1326_ (
  .in1({ S752, S744 }),
  .out1({ S754 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1327_ (
  .in1({ S753, S745 }),
  .out1({ S755 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1328_ (
  .in1({ S754, S731 }),
  .out1({ S756 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1329_ (
  .in1({ S755, S730 }),
  .out1({ S757 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1330_ (
  .in1({ S756, S726 }),
  .out1({ S758 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1331_ (
  .in1({ S757, S727 }),
  .out1({ S759 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1332_ (
  .in1({ S758, S717 }),
  .out1({ S760 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1333_ (
  .in1({ S759, S716 }),
  .out1({ S761 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1334_ (
  .in1({ S760, S712 }),
  .out1({ S762 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1335_ (
  .in1({ S761, S713 }),
  .out1({ S763 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1336_ (
  .in1({ S762, S705 }),
  .out1({ S764 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1337_ (
  .in1({ S763, S704 }),
  .out1({ S765 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1338_ (
  .in1({ S764, S700 }),
  .out1({ S766 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1339_ (
  .in1({ S765, S701 }),
  .out1({ S767 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1340_ (
  .in1({ S766, S693 }),
  .out1({ S768 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1341_ (
  .in1({ S767, S692 }),
  .out1({ S769 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1342_ (
  .in1({ S768, S688 }),
  .out1({ S770 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1343_ (
  .in1({ S769, S689 }),
  .out1({ S771 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1344_ (
  .in1({ S770, S678 }),
  .out1({ S772 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1345_ (
  .in1({ S771, S677 }),
  .out1({ S773 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1346_ (
  .in1({ S772, S673 }),
  .out1({ S774 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1347_ (
  .in1({ S773, S674 }),
  .out1({ S775 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1348_ (
  .in1({ S229, S222 }),
  .out1({ S776 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1349_ (
  .in1({ S775, S231 }),
  .out1({ S777 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1350_ (
  .in1({ S776, S774 }),
  .out1({ S778 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1351_ (
  .in1({ S778, S777 }),
  .out1({ S779 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1352_ (
  .in1({ S779, S654 }),
  .out1({ S780 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1353_ (
  .in1({ S547, S229 }),
  .out1({ S781 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1354_ (
  .in1({ S781, S222 }),
  .out1({ S782 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1355_ (
  .in1({ S782 }),
  .out1({ S783 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1356_ (
  .in1({ S782, S774 }),
  .out1({ S784 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1357_ (
  .in1({ S783, S775 }),
  .out1({ S785 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1358_ (
  .in1({ S653, S231 }),
  .out1({ S786 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1359_ (
  .in1({ S654, S230 }),
  .out1({ S787 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1360_ (
  .in1({ S786, S784 }),
  .out1({ S788 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1361_ (
  .in1({ S787, S785 }),
  .out1({ S789 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1362_ (
  .in1({ S770, S678 }),
  .out1({ S790 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1363_ (
  .in1({ S790, S773 }),
  .out1({ S791 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1364_ (
  .in1({ S791, S789 }),
  .out1({ S792 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1365_ (
  .in1({ S788, S672 }),
  .out1({ S793 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1366_ (
  .in1({ S793, S792 }),
  .out1({ S794 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1367_ (
  .in1({ S794 }),
  .out1({ S795 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1368_ (
  .in1({ S794, S229 }),
  .out1({ S796 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1369_ (
  .in1({ S795, S228 }),
  .out1({ S797 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1370_ (
  .in1({ S794, S229 }),
  .out1({ S798 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1371_ (
  .in1({ S798, S797 }),
  .out1({ S799 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1372_ (
  .in1({ S799 }),
  .out1({ S800 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1373_ (
  .in1({ S766, S693 }),
  .out1({ S801 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1374_ (
  .in1({ S801 }),
  .out1({ S802 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1375_ (
  .in1({ S802, S768 }),
  .out1({ S803 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1376_ (
  .in1({ S803, S788 }),
  .out1({ S804 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1377_ (
  .in1({ S804 }),
  .out1({ S805 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1378_ (
  .in1({ S789, S686 }),
  .out1({ S806 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1379_ (
  .in1({ S788, S687 }),
  .out1({ S807 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1380_ (
  .in1({ S806, S804 }),
  .out1({ S808 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1381_ (
  .in1({ S807, S805 }),
  .out1({ S809 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1382_ (
  .in1({ S809, S203 }),
  .out1({ S810 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1383_ (
  .in1({ S808, S202 }),
  .out1({ S811 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1384_ (
  .in1({ S808, S202 }),
  .out1({ S812 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1385_ (
  .in1({ S809, S203 }),
  .out1({ S813 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1386_ (
  .in1({ S763, S704 }),
  .out1({ S814 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1387_ (
  .in1({ S814, S764 }),
  .out1({ S815 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1388_ (
  .in1({ S815, S788 }),
  .out1({ S816 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1389_ (
  .in1({ S816 }),
  .out1({ S817 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1390_ (
  .in1({ S788, S698 }),
  .out1({ S818 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1391_ (
  .in1({ S818 }),
  .out1({ S819 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1392_ (
  .in1({ S819, S816 }),
  .out1({ S820 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1393_ (
  .in1({ S818, S817 }),
  .out1({ S821 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1394_ (
  .in1({ S821, S209 }),
  .out1({ S822 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1395_ (
  .in1({ S820, S208 }),
  .out1({ S823 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1396_ (
  .in1({ S820, S208 }),
  .out1({ S824 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1397_ (
  .in1({ S821, S209 }),
  .out1({ S825 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1398_ (
  .in1({ S824, S822 }),
  .out1({ S826 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1399_ (
  .in1({ S825, S823 }),
  .out1({ S827 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1400_ (
  .in1({ S759, S716 }),
  .out1({ S828 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1401_ (
  .in1({ S828, S760 }),
  .out1({ S829 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1402_ (
  .in1({ S829, S788 }),
  .out1({ S830 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1403_ (
  .in1({ S830 }),
  .out1({ S831 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1404_ (
  .in1({ S788, S710 }),
  .out1({ S832 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1405_ (
  .in1({ S832 }),
  .out1({ S833 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1406_ (
  .in1({ S833, S830 }),
  .out1({ S834 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1407_ (
  .in1({ S832, S831 }),
  .out1({ S835 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1408_ (
  .in1({ S835, S241 }),
  .out1({ S836 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1409_ (
  .in1({ S834, S240 }),
  .out1({ S837 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1410_ (
  .in1({ S834, S240 }),
  .out1({ S838 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1411_ (
  .in1({ S835, S241 }),
  .out1({ S839 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1412_ (
  .in1({ S838, S836 }),
  .out1({ S840 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1413_ (
  .in1({ S839, S837 }),
  .out1({ S841 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1414_ (
  .in1({ S755, S730 }),
  .out1({ S842 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1415_ (
  .in1({ S842, S756 }),
  .out1({ S843 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1416_ (
  .in1({ S843, S788 }),
  .out1({ S844 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1417_ (
  .in1({ S844 }),
  .out1({ S845 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1418_ (
  .in1({ S789, S724 }),
  .out1({ S846 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1419_ (
  .in1({ S788, S725 }),
  .out1({ S847 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1420_ (
  .in1({ S846, S844 }),
  .out1({ S848 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1421_ (
  .in1({ S847, S845 }),
  .out1({ S849 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1422_ (
  .in1({ S849, S249 }),
  .out1({ S850 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1423_ (
  .in1({ S848, S248 }),
  .out1({ S851 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1424_ (
  .in1({ S848, S248 }),
  .out1({ S852 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1425_ (
  .in1({ S849, S249 }),
  .out1({ S853 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1426_ (
  .in1({ S852, S850 }),
  .out1({ S854 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1427_ (
  .in1({ S853, S851 }),
  .out1({ S855 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1428_ (
  .in1({ S750, S747 }),
  .out1({ S856 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1429_ (
  .in1({ S856, S752 }),
  .out1({ S857 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1430_ (
  .in1({ S857, S788 }),
  .out1({ S858 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1431_ (
  .in1({ S858 }),
  .out1({ S859 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1432_ (
  .in1({ S789, S742 }),
  .out1({ S860 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1433_ (
  .in1({ S788, S743 }),
  .out1({ S861 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1434_ (
  .in1({ S860, S858 }),
  .out1({ S862 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1435_ (
  .in1({ S861, S859 }),
  .out1({ S863 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1436_ (
  .in1({ S863, S257 }),
  .out1({ S864 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1437_ (
  .in1({ S862, S256 }),
  .out1({ S865 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1438_ (
  .in1({ S862, S256 }),
  .out1({ S866 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1439_ (
  .in1({ S863, S257 }),
  .out1({ S867 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1440_ (
  .in1({ S271, S3325 }),
  .out1({ S868 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1441_ (
  .in1({ S270, new_datapath_addsubunit_in1_8 }),
  .out1({ S869 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1442_ (
  .in1({ S868, S746 }),
  .out1({ S870 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1443_ (
  .in1({ S869, S747 }),
  .out1({ S871 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1444_ (
  .in1({ S871, S788 }),
  .out1({ S872 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1445_ (
  .in1({ S870, S789 }),
  .out1({ S873 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1446_ (
  .in1({ S789, new_datapath_addsubunit_in1_8 }),
  .out1({ S874 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1447_ (
  .in1({ S788, S3325 }),
  .out1({ S875 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1448_ (
  .in1({ S874, S872 }),
  .out1({ S876 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1449_ (
  .in1({ S875, S873 }),
  .out1({ S877 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1450_ (
  .in1({ S877, S265 }),
  .out1({ S878 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1451_ (
  .in1({ S876, S264 }),
  .out1({ S879 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1452_ (
  .in1({ S270, new_datapath_addsubunit_in1_6 }),
  .out1({ S880 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1453_ (
  .in1({ S271, S5916 }),
  .out1({ S881 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1454_ (
  .in1({ S270, S5916 }),
  .out1({ S882 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1455_ (
  .in1({ S271, new_datapath_addsubunit_in1_6 }),
  .out1({ S883 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1456_ (
  .in1({ S271, new_datapath_addsubunit_in1_7 }),
  .out1({ S884 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1457_ (
  .in1({ S270, S5907 }),
  .out1({ S885 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1458_ (
  .in1({ S270, S5907 }),
  .out1({ S886 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1459_ (
  .in1({ S271, new_datapath_addsubunit_in1_7 }),
  .out1({ S887 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1460_ (
  .in1({ S886, S884 }),
  .out1({ S888 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1461_ (
  .in1({ S887, S885 }),
  .out1({ S889 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1462_ (
  .in1({ S270, new_datapath_addsubunit_in1_7 }),
  .out1({ S890 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1463_ (
  .in1({ S271, S5907 }),
  .out1({ S891 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1464_ (
  .in1({ S876, S264 }),
  .out1({ S892 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1465_ (
  .in1({ S877, S265 }),
  .out1({ S893 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1466_ (
  .in1({ S892, S878 }),
  .out1({ S894 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1467_ (
  .in1({ S893, S879 }),
  .out1({ S895 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1468_ (
  .in1({ S895, S890 }),
  .out1({ S896 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1469_ (
  .in1({ S894, S891 }),
  .out1({ S897 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1470_ (
  .in1({ S896, S878 }),
  .out1({ S898 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1471_ (
  .in1({ S897, S879 }),
  .out1({ S899 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1472_ (
  .in1({ S898, S866 }),
  .out1({ S900 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1473_ (
  .in1({ S899, S867 }),
  .out1({ S901 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1474_ (
  .in1({ S900, S864 }),
  .out1({ S902 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1475_ (
  .in1({ S901, S865 }),
  .out1({ S903 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1476_ (
  .in1({ S902, S855 }),
  .out1({ S904 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1477_ (
  .in1({ S903, S854 }),
  .out1({ S905 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1478_ (
  .in1({ S904, S850 }),
  .out1({ S906 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1479_ (
  .in1({ S905, S851 }),
  .out1({ S907 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1480_ (
  .in1({ S906, S841 }),
  .out1({ S908 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1481_ (
  .in1({ S907, S840 }),
  .out1({ S909 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1482_ (
  .in1({ S908, S836 }),
  .out1({ S910 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1483_ (
  .in1({ S909, S837 }),
  .out1({ S911 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1484_ (
  .in1({ S910, S827 }),
  .out1({ S912 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1485_ (
  .in1({ S911, S826 }),
  .out1({ S913 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1486_ (
  .in1({ S912, S822 }),
  .out1({ S914 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1487_ (
  .in1({ S913, S823 }),
  .out1({ S915 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1488_ (
  .in1({ S914, S812 }),
  .out1({ S916 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1489_ (
  .in1({ S915, S813 }),
  .out1({ S917 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1490_ (
  .in1({ S916, S810 }),
  .out1({ S918 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1491_ (
  .in1({ S917, S811 }),
  .out1({ S919 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1492_ (
  .in1({ S918, S799 }),
  .out1({ S920 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1493_ (
  .in1({ S919, S800 }),
  .out1({ S921 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1494_ (
  .in1({ S920, S796 }),
  .out1({ S922 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1495_ (
  .in1({ S921, S797 }),
  .out1({ S923 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1496_ (
  .in1({ S220, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S924 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1497_ (
  .in1({ S922, S222 }),
  .out1({ S925 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1498_ (
  .in1({ S924, S922 }),
  .out1({ S926 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1499_ (
  .in1({ S926, S780 }),
  .out1({ S927 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1500_ (
  .in1({ S927, S925 }),
  .out1({ S928 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1501_ (
  .in1({ S780, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S929 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1502_ (
  .in1({ S929 }),
  .out1({ S930 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1503_ (
  .in1({ S929, S923 }),
  .out1({ S931 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1504_ (
  .in1({ S930, S922 }),
  .out1({ S932 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1505_ (
  .in1({ S653, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S933 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1506_ (
  .in1({ S933, S220 }),
  .out1({ S934 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1507_ (
  .in1({ S934 }),
  .out1({ S935 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1508_ (
  .in1({ S934, S931 }),
  .out1({ S936 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1509_ (
  .in1({ S935, S932 }),
  .out1({ S937 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1510_ (
  .in1({ S918, S799 }),
  .out1({ S938 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1511_ (
  .in1({ S938, S921 }),
  .out1({ S939 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1512_ (
  .in1({ S939, S936 }),
  .out1({ S940 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1513_ (
  .in1({ S937, S794 }),
  .out1({ S941 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1514_ (
  .in1({ S941, S940 }),
  .out1({ S942 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1515_ (
  .in1({ S942 }),
  .out1({ S943 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1516_ (
  .in1({ S942, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S944 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1517_ (
  .in1({ S943, S3478 }),
  .out1({ S945 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1518_ (
  .in1({ S942, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S946 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1519_ (
  .in1({ S946 }),
  .out1({ S947 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1520_ (
  .in1({ S947, S944 }),
  .out1({ S948 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1521_ (
  .in1({ S948 }),
  .out1({ S949 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1522_ (
  .in1({ S812, S810 }),
  .out1({ S950 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1523_ (
  .in1({ S813, S811 }),
  .out1({ S951 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1524_ (
  .in1({ S951, S914 }),
  .out1({ S952 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1525_ (
  .in1({ S950, S915 }),
  .out1({ S953 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1526_ (
  .in1({ S953, S952 }),
  .out1({ S954 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1527_ (
  .in1({ S954, S936 }),
  .out1({ S955 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1528_ (
  .in1({ S937, S809 }),
  .out1({ S956 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1529_ (
  .in1({ S956, S955 }),
  .out1({ S957 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1530_ (
  .in1({ S957 }),
  .out1({ S958 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1531_ (
  .in1({ S957, S229 }),
  .out1({ S959 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1532_ (
  .in1({ S958, S228 }),
  .out1({ S960 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1533_ (
  .in1({ S958, S228 }),
  .out1({ S961 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1534_ (
  .in1({ S957, S229 }),
  .out1({ S962 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1535_ (
  .in1({ S911, S826 }),
  .out1({ S963 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1536_ (
  .in1({ S963, S912 }),
  .out1({ S964 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1537_ (
  .in1({ S964, S937 }),
  .out1({ S965 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1538_ (
  .in1({ S965 }),
  .out1({ S966 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1539_ (
  .in1({ S937, S821 }),
  .out1({ S967 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1540_ (
  .in1({ S967 }),
  .out1({ S968 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1541_ (
  .in1({ S968, S965 }),
  .out1({ S969 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1542_ (
  .in1({ S967, S966 }),
  .out1({ S970 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1543_ (
  .in1({ S970, S203 }),
  .out1({ S971 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1544_ (
  .in1({ S969, S202 }),
  .out1({ S972 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1545_ (
  .in1({ S969, S202 }),
  .out1({ S973 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1546_ (
  .in1({ S970, S203 }),
  .out1({ S974 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1547_ (
  .in1({ S973, S971 }),
  .out1({ S975 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1548_ (
  .in1({ S974, S972 }),
  .out1({ S976 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1549_ (
  .in1({ S906, S841 }),
  .out1({ S977 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1550_ (
  .in1({ S977, S909 }),
  .out1({ S978 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1551_ (
  .in1({ S978, S936 }),
  .out1({ S979 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1552_ (
  .in1({ S937, S835 }),
  .out1({ S980 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1553_ (
  .in1({ S980, S979 }),
  .out1({ S981 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1554_ (
  .in1({ S981 }),
  .out1({ S982 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1555_ (
  .in1({ S981, S209 }),
  .out1({ S983 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1556_ (
  .in1({ S982, S208 }),
  .out1({ S984 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1557_ (
  .in1({ S982, S208 }),
  .out1({ S985 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1558_ (
  .in1({ S985, S983 }),
  .out1({ S986 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1559_ (
  .in1({ S986 }),
  .out1({ S987 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1560_ (
  .in1({ S903, S854 }),
  .out1({ S988 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1561_ (
  .in1({ S988, S904 }),
  .out1({ S989 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1562_ (
  .in1({ S989, S937 }),
  .out1({ S990 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1563_ (
  .in1({ S990 }),
  .out1({ S991 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1564_ (
  .in1({ S936, S848 }),
  .out1({ S992 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1565_ (
  .in1({ S937, S849 }),
  .out1({ S993 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1566_ (
  .in1({ S992, S990 }),
  .out1({ S994 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1567_ (
  .in1({ S993, S991 }),
  .out1({ S995 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1568_ (
  .in1({ S995, S241 }),
  .out1({ S996 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1569_ (
  .in1({ S994, S240 }),
  .out1({ S997 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1570_ (
  .in1({ S994, S240 }),
  .out1({ S998 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1571_ (
  .in1({ S995, S241 }),
  .out1({ S999 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1572_ (
  .in1({ S998, S996 }),
  .out1({ S1000 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1573_ (
  .in1({ S999, S997 }),
  .out1({ S1001 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1574_ (
  .in1({ S866, S864 }),
  .out1({ S1002 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1575_ (
  .in1({ S867, S865 }),
  .out1({ S1003 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1576_ (
  .in1({ S1002, S898 }),
  .out1({ S1004 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1577_ (
  .in1({ S1003, S899 }),
  .out1({ S1005 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1578_ (
  .in1({ S1005, S1004 }),
  .out1({ S1006 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1579_ (
  .in1({ S1006, S937 }),
  .out1({ S1007 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1580_ (
  .in1({ S1007 }),
  .out1({ S1008 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1581_ (
  .in1({ S936, S862 }),
  .out1({ S1009 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1582_ (
  .in1({ S937, S863 }),
  .out1({ S1010 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1583_ (
  .in1({ S1009, S1007 }),
  .out1({ S1011 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1584_ (
  .in1({ S1010, S1008 }),
  .out1({ S1012 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1585_ (
  .in1({ S1012, S249 }),
  .out1({ S1013 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1586_ (
  .in1({ S1011, S248 }),
  .out1({ S1014 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1587_ (
  .in1({ S894, S891 }),
  .out1({ S1015 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1588_ (
  .in1({ S1015, S896 }),
  .out1({ S1016 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1589_ (
  .in1({ S1016, S937 }),
  .out1({ S1017 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1590_ (
  .in1({ S1017 }),
  .out1({ S1018 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1591_ (
  .in1({ S936, S876 }),
  .out1({ S1019 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1592_ (
  .in1({ S937, S877 }),
  .out1({ S1020 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1593_ (
  .in1({ S1019, S1017 }),
  .out1({ S1021 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1594_ (
  .in1({ S1020, S1018 }),
  .out1({ S1022 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1595_ (
  .in1({ S1022, S257 }),
  .out1({ S1023 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1596_ (
  .in1({ S1021, S256 }),
  .out1({ S1024 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1597_ (
  .in1({ S937, S889 }),
  .out1({ S1025 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1598_ (
  .in1({ S936, S888 }),
  .out1({ S1026 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1599_ (
  .in1({ S936, S5907 }),
  .out1({ S1027 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1600_ (
  .in1({ S937, new_datapath_addsubunit_in1_7 }),
  .out1({ S1028 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1601_ (
  .in1({ S1027, S1025 }),
  .out1({ S1029 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1602_ (
  .in1({ S1028, S1026 }),
  .out1({ S1030 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1603_ (
  .in1({ S1029, S265 }),
  .out1({ S1031 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1604_ (
  .in1({ S1030, S264 }),
  .out1({ S1032 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1605_ (
  .in1({ S1030, S264 }),
  .out1({ S1033 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1606_ (
  .in1({ S1029, S265 }),
  .out1({ S1034 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1607_ (
  .in1({ S1033, S1031 }),
  .out1({ S1035 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1608_ (
  .in1({ S1034, S1032 }),
  .out1({ S1036 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1609_ (
  .in1({ S1036, S880 }),
  .out1({ S1037 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1610_ (
  .in1({ S1035, S881 }),
  .out1({ S1038 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1611_ (
  .in1({ S1037, S1031 }),
  .out1({ S1039 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1612_ (
  .in1({ S1038, S1032 }),
  .out1({ S1040 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1613_ (
  .in1({ S1021, S256 }),
  .out1({ S1041 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1614_ (
  .in1({ S1041, S1023 }),
  .out1({ S1042 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1615_ (
  .in1({ S1042 }),
  .out1({ S1043 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1616_ (
  .in1({ S1043, S1039 }),
  .out1({ S1044 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1617_ (
  .in1({ S1042, S1040 }),
  .out1({ S1045 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1618_ (
  .in1({ S1044, S1023 }),
  .out1({ S1046 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1619_ (
  .in1({ S1045, S1024 }),
  .out1({ S1047 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1620_ (
  .in1({ S1046, S1014 }),
  .out1({ S1048 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1621_ (
  .in1({ S1047, S1013 }),
  .out1({ S1049 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1622_ (
  .in1({ S1048, S1013 }),
  .out1({ S1050 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1623_ (
  .in1({ S1049, S1014 }),
  .out1({ S1051 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1624_ (
  .in1({ S1050, S1001 }),
  .out1({ S1052 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1625_ (
  .in1({ S1051, S1000 }),
  .out1({ S1053 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1626_ (
  .in1({ S1052, S996 }),
  .out1({ S1054 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1627_ (
  .in1({ S1053, S997 }),
  .out1({ S1055 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1628_ (
  .in1({ S1054, S987 }),
  .out1({ S1056 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1629_ (
  .in1({ S1055, S986 }),
  .out1({ S1057 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1630_ (
  .in1({ S1056, S983 }),
  .out1({ S1058 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1631_ (
  .in1({ S1057, S984 }),
  .out1({ S1059 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1632_ (
  .in1({ S1058, S976 }),
  .out1({ S1060 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1633_ (
  .in1({ S1059, S975 }),
  .out1({ S1061 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1634_ (
  .in1({ S1060, S971 }),
  .out1({ S1062 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1635_ (
  .in1({ S1061, S972 }),
  .out1({ S1063 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1636_ (
  .in1({ S1062, S961 }),
  .out1({ S1064 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1637_ (
  .in1({ S1063, S962 }),
  .out1({ S1065 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1638_ (
  .in1({ S1064, S959 }),
  .out1({ S1066 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1639_ (
  .in1({ S1065, S960 }),
  .out1({ S1067 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1640_ (
  .in1({ S1066, S949 }),
  .out1({ S1068 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1641_ (
  .in1({ S1067, S948 }),
  .out1({ S1069 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1642_ (
  .in1({ S1068, S944 }),
  .out1({ S1070 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1643_ (
  .in1({ S1069, S945 }),
  .out1({ S1071 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1644_ (
  .in1({ S218, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S1072 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1645_ (
  .in1({ S1070, S220 }),
  .out1({ S1073 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1646_ (
  .in1({ S1072, S1070 }),
  .out1({ S1074 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1647_ (
  .in1({ S1074, S928 }),
  .out1({ S1075 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1648_ (
  .in1({ S1075, S1073 }),
  .out1({ S1076 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1649_ (
  .in1({ S928, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S1077 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1650_ (
  .in1({ S1077 }),
  .out1({ S1078 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1651_ (
  .in1({ S1077, S1071 }),
  .out1({ S1079 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1652_ (
  .in1({ S1078, S1070 }),
  .out1({ S1080 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1653_ (
  .in1({ S780, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S1081 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1654_ (
  .in1({ S1081, S218 }),
  .out1({ S1082 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1655_ (
  .in1({ S1082 }),
  .out1({ S1083 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1656_ (
  .in1({ S1082, S1079 }),
  .out1({ S1084 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1657_ (
  .in1({ S1083, S1080 }),
  .out1({ S1085 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1658_ (
  .in1({ S1066, S949 }),
  .out1({ S1086 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1659_ (
  .in1({ S1086, S1069 }),
  .out1({ S1087 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1660_ (
  .in1({ S1087, S1084 }),
  .out1({ S1088 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1661_ (
  .in1({ S1085, S942 }),
  .out1({ S1089 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1662_ (
  .in1({ S1089, S1088 }),
  .out1({ S1090 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1663_ (
  .in1({ S1090 }),
  .out1({ S1091 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1664_ (
  .in1({ S1090, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S1092 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1665_ (
  .in1({ S1091, S3467 }),
  .out1({ S1093 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1666_ (
  .in1({ S1090, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S1094 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1667_ (
  .in1({ S1094, S1093 }),
  .out1({ S1095 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1668_ (
  .in1({ S1095 }),
  .out1({ S1096 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1669_ (
  .in1({ S961, S959 }),
  .out1({ S1097 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1670_ (
  .in1({ S962, S960 }),
  .out1({ S1098 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1671_ (
  .in1({ S1097, S1063 }),
  .out1({ S1099 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1672_ (
  .in1({ S1098, S1062 }),
  .out1({ S1100 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1673_ (
  .in1({ S1100, S1099 }),
  .out1({ S1101 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1674_ (
  .in1({ S1101, S1085 }),
  .out1({ S1102 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1675_ (
  .in1({ S1102 }),
  .out1({ S1103 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1676_ (
  .in1({ S1085, S957 }),
  .out1({ S1104 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1677_ (
  .in1({ S1104 }),
  .out1({ S1105 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1678_ (
  .in1({ S1105, S1102 }),
  .out1({ S1106 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1679_ (
  .in1({ S1104, S1103 }),
  .out1({ S1107 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1680_ (
  .in1({ S1107, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S1108 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1681_ (
  .in1({ S1106, S3478 }),
  .out1({ S1109 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1682_ (
  .in1({ S1058, S976 }),
  .out1({ S1110 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1683_ (
  .in1({ S1110, S1061 }),
  .out1({ S1111 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1684_ (
  .in1({ S1111, S1084 }),
  .out1({ S1112 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1685_ (
  .in1({ S1085, S970 }),
  .out1({ S1113 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1686_ (
  .in1({ S1113, S1112 }),
  .out1({ S1114 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1687_ (
  .in1({ S1114 }),
  .out1({ S1115 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1688_ (
  .in1({ S1114, S229 }),
  .out1({ S1116 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1689_ (
  .in1({ S1115, S228 }),
  .out1({ S1117 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1690_ (
  .in1({ S1114, S229 }),
  .out1({ S1118 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1691_ (
  .in1({ S1118, S1117 }),
  .out1({ S1119 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1692_ (
  .in1({ S1119 }),
  .out1({ S1120 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1693_ (
  .in1({ S1055, S986 }),
  .out1({ S1121 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1694_ (
  .in1({ S1121, S1056 }),
  .out1({ S1122 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1695_ (
  .in1({ S1122, S1085 }),
  .out1({ S1123 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1696_ (
  .in1({ S1123 }),
  .out1({ S1124 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1697_ (
  .in1({ S1085, S981 }),
  .out1({ S1125 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1698_ (
  .in1({ S1125 }),
  .out1({ S1126 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1699_ (
  .in1({ S1126, S1123 }),
  .out1({ S1127 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1700_ (
  .in1({ S1125, S1124 }),
  .out1({ S1128 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1701_ (
  .in1({ S1128, S203 }),
  .out1({ S1129 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1702_ (
  .in1({ S1127, S202 }),
  .out1({ S1130 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1703_ (
  .in1({ S1127, S202 }),
  .out1({ S1131 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1704_ (
  .in1({ S1128, S203 }),
  .out1({ S1132 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1705_ (
  .in1({ S1131, S1129 }),
  .out1({ S1133 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1706_ (
  .in1({ S1132, S1130 }),
  .out1({ S1134 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1707_ (
  .in1({ S1051, S1000 }),
  .out1({ S1135 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1708_ (
  .in1({ S1135, S1052 }),
  .out1({ S1136 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1709_ (
  .in1({ S1136, S1085 }),
  .out1({ S1137 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1710_ (
  .in1({ S1137 }),
  .out1({ S1138 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1711_ (
  .in1({ S1084, S994 }),
  .out1({ S1139 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1712_ (
  .in1({ S1085, S995 }),
  .out1({ S1140 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1713_ (
  .in1({ S1139, S1137 }),
  .out1({ S1141 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1714_ (
  .in1({ S1140, S1138 }),
  .out1({ S1142 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1715_ (
  .in1({ S1142, S209 }),
  .out1({ S1143 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1716_ (
  .in1({ S1141, S208 }),
  .out1({ S1144 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1717_ (
  .in1({ S1141, S208 }),
  .out1({ S1145 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1718_ (
  .in1({ S1142, S209 }),
  .out1({ S1146 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1719_ (
  .in1({ S1145, S1143 }),
  .out1({ S1147 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1720_ (
  .in1({ S1146, S1144 }),
  .out1({ S1148 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1721_ (
  .in1({ S1014, S1013 }),
  .out1({ S1149 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1722_ (
  .in1({ S1149, S1046 }),
  .out1({ S1150 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1723_ (
  .in1({ S1149, S1046 }),
  .out1({ S1151 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1724_ (
  .in1({ S1151 }),
  .out1({ S1152 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1725_ (
  .in1({ S1152, S1150 }),
  .out1({ S1153 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1726_ (
  .in1({ S1153, S1085 }),
  .out1({ S1154 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1727_ (
  .in1({ S1154 }),
  .out1({ S1155 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1728_ (
  .in1({ S1084, S1011 }),
  .out1({ S1156 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1729_ (
  .in1({ S1085, S1012 }),
  .out1({ S1157 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1730_ (
  .in1({ S1156, S1154 }),
  .out1({ S1158 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1731_ (
  .in1({ S1157, S1155 }),
  .out1({ S1159 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1732_ (
  .in1({ S1159, S241 }),
  .out1({ S1160 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1733_ (
  .in1({ S1158, S240 }),
  .out1({ S1161 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1734_ (
  .in1({ S1158, S240 }),
  .out1({ S1162 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1735_ (
  .in1({ S1159, S241 }),
  .out1({ S1163 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1736_ (
  .in1({ S1162, S1160 }),
  .out1({ S1164 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1737_ (
  .in1({ S1163, S1161 }),
  .out1({ S1165 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1738_ (
  .in1({ S1042, S1040 }),
  .out1({ S1166 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1739_ (
  .in1({ S1166, S1044 }),
  .out1({ S1167 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1740_ (
  .in1({ S1167, S1085 }),
  .out1({ S1168 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1741_ (
  .in1({ S1168 }),
  .out1({ S1169 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1742_ (
  .in1({ S1085, S1022 }),
  .out1({ S1170 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1743_ (
  .in1({ S1170 }),
  .out1({ S1171 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1744_ (
  .in1({ S1171, S1168 }),
  .out1({ S1172 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1745_ (
  .in1({ S1170, S1169 }),
  .out1({ S1173 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1746_ (
  .in1({ S1173, S249 }),
  .out1({ S1174 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1747_ (
  .in1({ S1172, S248 }),
  .out1({ S1175 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1748_ (
  .in1({ S1035, S881 }),
  .out1({ S1176 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1749_ (
  .in1({ S1176, S1037 }),
  .out1({ S1177 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1750_ (
  .in1({ S1177, S1085 }),
  .out1({ S1178 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1751_ (
  .in1({ S1084, S1030 }),
  .out1({ S1179 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1752_ (
  .in1({ S1179, S1178 }),
  .out1({ S1180 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1753_ (
  .in1({ S1180 }),
  .out1({ S1181 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1754_ (
  .in1({ S1181, S257 }),
  .out1({ S1182 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1755_ (
  .in1({ S1180, S256 }),
  .out1({ S1183 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1756_ (
  .in1({ S1180, S256 }),
  .out1({ S1184 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1757_ (
  .in1({ S1181, S257 }),
  .out1({ S1185 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1758_ (
  .in1({ S1184, S1182 }),
  .out1({ S1186 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1759_ (
  .in1({ S1185, S1183 }),
  .out1({ S1187 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1760_ (
  .in1({ S1085, S270 }),
  .out1({ S1188 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1761_ (
  .in1({ S1084, S271 }),
  .out1({ S1189 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1762_ (
  .in1({ S1188, S5916 }),
  .out1({ S1190 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1763_ (
  .in1({ S1189, new_datapath_addsubunit_in1_6 }),
  .out1({ S1191 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1764_ (
  .in1({ S1085, S881 }),
  .out1({ S1192 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1765_ (
  .in1({ S1084, S880 }),
  .out1({ S1193 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1766_ (
  .in1({ S1192, S1190 }),
  .out1({ S1194 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1767_ (
  .in1({ S1193, S1191 }),
  .out1({ S1195 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1768_ (
  .in1({ S1194, S265 }),
  .out1({ S1196 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1769_ (
  .in1({ S1195, S264 }),
  .out1({ S1197 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1770_ (
  .in1({ S1195, S264 }),
  .out1({ S1198 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1771_ (
  .in1({ S1194, S265 }),
  .out1({ S1199 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1772_ (
  .in1({ S1198, S1196 }),
  .out1({ S1200 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1773_ (
  .in1({ S1199, S1197 }),
  .out1({ S1201 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1774_ (
  .in1({ S270, new_datapath_addsubunit_in1_4 }),
  .out1({ S1202 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1775_ (
  .in1({ S271, S5936 }),
  .out1({ S1203 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1776_ (
  .in1({ S270, S5936 }),
  .out1({ S1204 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1777_ (
  .in1({ S271, new_datapath_addsubunit_in1_4 }),
  .out1({ S1205 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1778_ (
  .in1({ S271, new_datapath_addsubunit_in1_5 }),
  .out1({ S1206 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1779_ (
  .in1({ S270, S5926 }),
  .out1({ S1207 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1780_ (
  .in1({ S270, S5926 }),
  .out1({ S1208 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1781_ (
  .in1({ S271, new_datapath_addsubunit_in1_5 }),
  .out1({ S1209 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1782_ (
  .in1({ S1208, S1206 }),
  .out1({ S1210 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1783_ (
  .in1({ S1209, S1207 }),
  .out1({ S1211 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1784_ (
  .in1({ S270, new_datapath_addsubunit_in1_5 }),
  .out1({ S1212 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1785_ (
  .in1({ S271, S5926 }),
  .out1({ S1213 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1786_ (
  .in1({ S1212, S1201 }),
  .out1({ S1214 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1787_ (
  .in1({ S1213, S1200 }),
  .out1({ S1215 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1788_ (
  .in1({ S1214, S1196 }),
  .out1({ S1216 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1789_ (
  .in1({ S1215, S1197 }),
  .out1({ S1217 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1790_ (
  .in1({ S1216, S1187 }),
  .out1({ S1218 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1791_ (
  .in1({ S1217, S1186 }),
  .out1({ S1219 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1792_ (
  .in1({ S1218, S1182 }),
  .out1({ S1220 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1793_ (
  .in1({ S1219, S1183 }),
  .out1({ S1221 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1794_ (
  .in1({ S1172, S248 }),
  .out1({ S1222 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1795_ (
  .in1({ S1173, S249 }),
  .out1({ S1223 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1796_ (
  .in1({ S1222, S1174 }),
  .out1({ S1224 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1797_ (
  .in1({ S1223, S1175 }),
  .out1({ S1225 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1798_ (
  .in1({ S1225, S1220 }),
  .out1({ S1226 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1799_ (
  .in1({ S1224, S1221 }),
  .out1({ S1227 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1800_ (
  .in1({ S1226, S1174 }),
  .out1({ S1228 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1801_ (
  .in1({ S1227, S1175 }),
  .out1({ S1229 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1802_ (
  .in1({ S1228, S1165 }),
  .out1({ S1230 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1803_ (
  .in1({ S1229, S1164 }),
  .out1({ S1231 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1804_ (
  .in1({ S1230, S1160 }),
  .out1({ S1232 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1805_ (
  .in1({ S1231, S1161 }),
  .out1({ S1233 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1806_ (
  .in1({ S1232, S1148 }),
  .out1({ S1234 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1807_ (
  .in1({ S1233, S1147 }),
  .out1({ S1235 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1808_ (
  .in1({ S1234, S1143 }),
  .out1({ S1236 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1809_ (
  .in1({ S1235, S1144 }),
  .out1({ S1237 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1810_ (
  .in1({ S1236, S1134 }),
  .out1({ S1238 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1811_ (
  .in1({ S1237, S1133 }),
  .out1({ S1239 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1812_ (
  .in1({ S1238, S1129 }),
  .out1({ S1240 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1813_ (
  .in1({ S1239, S1130 }),
  .out1({ S1241 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1814_ (
  .in1({ S1240, S1119 }),
  .out1({ S1242 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1815_ (
  .in1({ S1241, S1120 }),
  .out1({ S1243 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1816_ (
  .in1({ S1242, S1116 }),
  .out1({ S1244 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1817_ (
  .in1({ S1243, S1117 }),
  .out1({ S1245 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1818_ (
  .in1({ S1244, S1109 }),
  .out1({ S1246 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1819_ (
  .in1({ S1245, S1108 }),
  .out1({ S1247 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1820_ (
  .in1({ S1246, S1108 }),
  .out1({ S1248 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1821_ (
  .in1({ S1247, S1109 }),
  .out1({ S1249 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1822_ (
  .in1({ S1248, S1095 }),
  .out1({ S1250 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1823_ (
  .in1({ S1249, S1096 }),
  .out1({ S1251 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1824_ (
  .in1({ S1250, S1092 }),
  .out1({ S1252 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1825_ (
  .in1({ S1251, S1093 }),
  .out1({ S1253 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1826_ (
  .in1({ S216, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S1254 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1827_ (
  .in1({ S1252, S218 }),
  .out1({ S1255 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1828_ (
  .in1({ S1254, S1252 }),
  .out1({ S1256 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1829_ (
  .in1({ S1256, S1076 }),
  .out1({ S1257 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1830_ (
  .in1({ S1257, S1255 }),
  .out1({ S1258 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1831_ (
  .in1({ S1258 }),
  .out1({ S1259 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1832_ (
  .in1({ S1076, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S1260 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1833_ (
  .in1({ S1260 }),
  .out1({ S1261 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1834_ (
  .in1({ S1260, S1253 }),
  .out1({ S1262 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1835_ (
  .in1({ S1261, S1252 }),
  .out1({ S1263 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1836_ (
  .in1({ S928, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S1264 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1837_ (
  .in1({ S1264, S216 }),
  .out1({ S1265 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1838_ (
  .in1({ S1265 }),
  .out1({ S1266 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1839_ (
  .in1({ S1265, S1262 }),
  .out1({ S1267 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1840_ (
  .in1({ S1266, S1263 }),
  .out1({ S1268 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1841_ (
  .in1({ S1248, S1095 }),
  .out1({ S1269 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1842_ (
  .in1({ S1269, S1251 }),
  .out1({ S1270 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1843_ (
  .in1({ S1270, S1267 }),
  .out1({ S1271 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1844_ (
  .in1({ S1268, S1090 }),
  .out1({ S1272 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1845_ (
  .in1({ S1272, S1271 }),
  .out1({ S1273 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1846_ (
  .in1({ S1273 }),
  .out1({ S1274 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1847_ (
  .in1({ S1273, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S1275 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1848_ (
  .in1({ S1274, S3456 }),
  .out1({ S1276 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1849_ (
  .in1({ S1273, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S1277 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1850_ (
  .in1({ S1277, S1276 }),
  .out1({ S1278 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1851_ (
  .in1({ S1278 }),
  .out1({ S1279 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1852_ (
  .in1({ S1109, S1108 }),
  .out1({ S1280 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1853_ (
  .in1({ S1280, S1245 }),
  .out1({ S1281 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1854_ (
  .in1({ S1280, S1245 }),
  .out1({ S1282 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1855_ (
  .in1({ S1282 }),
  .out1({ S1283 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1856_ (
  .in1({ S1283, S1281 }),
  .out1({ S1284 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1857_ (
  .in1({ S1284, S1268 }),
  .out1({ S1285 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1858_ (
  .in1({ S1285 }),
  .out1({ S1286 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1859_ (
  .in1({ S1268, S1107 }),
  .out1({ S1287 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1860_ (
  .in1({ S1287 }),
  .out1({ S1288 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1861_ (
  .in1({ S1288, S1285 }),
  .out1({ S1289 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1862_ (
  .in1({ S1287, S1286 }),
  .out1({ S1290 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1863_ (
  .in1({ S1289, S3467 }),
  .out1({ S1291 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1864_ (
  .in1({ S1290, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S1292 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1865_ (
  .in1({ S1240, S1119 }),
  .out1({ S1293 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1866_ (
  .in1({ S1293, S1243 }),
  .out1({ S1294 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1867_ (
  .in1({ S1294, S1267 }),
  .out1({ S1295 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1868_ (
  .in1({ S1268, S1114 }),
  .out1({ S1296 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1869_ (
  .in1({ S1296, S1295 }),
  .out1({ S1297 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1870_ (
  .in1({ S1297 }),
  .out1({ S1298 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1871_ (
  .in1({ S1297, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S1299 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1872_ (
  .in1({ S1298, S3478 }),
  .out1({ S1300 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1873_ (
  .in1({ S1297, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S1301 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1874_ (
  .in1({ S1301, S1300 }),
  .out1({ S1302 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1875_ (
  .in1({ S1302 }),
  .out1({ S1303 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1876_ (
  .in1({ S1237, S1133 }),
  .out1({ S1304 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1877_ (
  .in1({ S1304, S1238 }),
  .out1({ S1305 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1878_ (
  .in1({ S1305, S1268 }),
  .out1({ S1306 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1879_ (
  .in1({ S1306 }),
  .out1({ S1307 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1880_ (
  .in1({ S1268, S1128 }),
  .out1({ S1308 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1881_ (
  .in1({ S1308 }),
  .out1({ S1309 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1882_ (
  .in1({ S1309, S1306 }),
  .out1({ S1310 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1883_ (
  .in1({ S1308, S1307 }),
  .out1({ S1311 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1884_ (
  .in1({ S1311, S229 }),
  .out1({ S1312 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1885_ (
  .in1({ S1310, S228 }),
  .out1({ S1313 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1886_ (
  .in1({ S1310, S228 }),
  .out1({ S1314 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1887_ (
  .in1({ S1311, S229 }),
  .out1({ S1315 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1888_ (
  .in1({ S1233, S1147 }),
  .out1({ S1316 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1889_ (
  .in1({ S1316, S1234 }),
  .out1({ S1317 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1890_ (
  .in1({ S1317, S1268 }),
  .out1({ S1318 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1891_ (
  .in1({ S1318 }),
  .out1({ S1319 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1892_ (
  .in1({ S1267, S1141 }),
  .out1({ S1320 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1893_ (
  .in1({ S1268, S1142 }),
  .out1({ S1321 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1894_ (
  .in1({ S1320, S1318 }),
  .out1({ S1322 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1895_ (
  .in1({ S1321, S1319 }),
  .out1({ S1323 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1896_ (
  .in1({ S1323, S203 }),
  .out1({ S1324 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1897_ (
  .in1({ S1322, S202 }),
  .out1({ S1325 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1898_ (
  .in1({ S1322, S202 }),
  .out1({ S1326 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1899_ (
  .in1({ S1323, S203 }),
  .out1({ S1327 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1900_ (
  .in1({ S1326, S1324 }),
  .out1({ S1328 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1901_ (
  .in1({ S1327, S1325 }),
  .out1({ S1329 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1902_ (
  .in1({ S1267, S1158 }),
  .out1({ S1330 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1903_ (
  .in1({ S1268, S1159 }),
  .out1({ S1331 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1904_ (
  .in1({ S1229, S1164 }),
  .out1({ S1332 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1905_ (
  .in1({ S1332, S1230 }),
  .out1({ S1333 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1906_ (
  .in1({ S1333, S1268 }),
  .out1({ S1334 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1907_ (
  .in1({ S1334 }),
  .out1({ S1335 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1908_ (
  .in1({ S1334, S1330 }),
  .out1({ S1336 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1909_ (
  .in1({ S1335, S1331 }),
  .out1({ S1337 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1910_ (
  .in1({ S1337, S209 }),
  .out1({ S1338 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1911_ (
  .in1({ S1336, S208 }),
  .out1({ S1339 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1912_ (
  .in1({ S1336, S208 }),
  .out1({ S1340 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1913_ (
  .in1({ S1337, S209 }),
  .out1({ S1341 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1914_ (
  .in1({ S1340, S1338 }),
  .out1({ S1342 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1915_ (
  .in1({ S1341, S1339 }),
  .out1({ S1343 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1916_ (
  .in1({ S1268, S1173 }),
  .out1({ S1344 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1917_ (
  .in1({ S1344 }),
  .out1({ S1345 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1918_ (
  .in1({ S1224, S1221 }),
  .out1({ S1346 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1919_ (
  .in1({ S1346, S1226 }),
  .out1({ S1347 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1920_ (
  .in1({ S1347, S1268 }),
  .out1({ S1348 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1921_ (
  .in1({ S1348 }),
  .out1({ S1349 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1922_ (
  .in1({ S1348, S1345 }),
  .out1({ S1350 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1923_ (
  .in1({ S1349, S1344 }),
  .out1({ S1351 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1924_ (
  .in1({ S1351, S241 }),
  .out1({ S1352 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1925_ (
  .in1({ S1350, S240 }),
  .out1({ S1353 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1926_ (
  .in1({ S1267, S1180 }),
  .out1({ S1354 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1927_ (
  .in1({ S1268, S1181 }),
  .out1({ S1355 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1928_ (
  .in1({ S1217, S1186 }),
  .out1({ S1356 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1929_ (
  .in1({ S1356, S1218 }),
  .out1({ S1357 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1930_ (
  .in1({ S1357, S1268 }),
  .out1({ S1358 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1931_ (
  .in1({ S1358 }),
  .out1({ S1359 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1932_ (
  .in1({ S1358, S1354 }),
  .out1({ S1360 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1933_ (
  .in1({ S1359, S1355 }),
  .out1({ S1361 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1934_ (
  .in1({ S1361, S249 }),
  .out1({ S1362 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1935_ (
  .in1({ S1360, S248 }),
  .out1({ S1363 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1936_ (
  .in1({ S1360, S248 }),
  .out1({ S1364 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1937_ (
  .in1({ S1361, S249 }),
  .out1({ S1365 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1938_ (
  .in1({ S1364, S1362 }),
  .out1({ S1366 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1939_ (
  .in1({ S1365, S1363 }),
  .out1({ S1367 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1940_ (
  .in1({ S1213, S1200 }),
  .out1({ S1368 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1941_ (
  .in1({ S1368, S1214 }),
  .out1({ S1369 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1942_ (
  .in1({ S1369, S1268 }),
  .out1({ S1370 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1943_ (
  .in1({ S1370 }),
  .out1({ S1371 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1944_ (
  .in1({ S1268, S1194 }),
  .out1({ S1372 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_1945_ (
  .in1({ S1372 }),
  .out1({ S1373 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1946_ (
  .in1({ S1373, S1370 }),
  .out1({ S1374 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1947_ (
  .in1({ S1372, S1371 }),
  .out1({ S1375 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1948_ (
  .in1({ S1375, S257 }),
  .out1({ S1376 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1949_ (
  .in1({ S1374, S256 }),
  .out1({ S1377 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1950_ (
  .in1({ S1374, S256 }),
  .out1({ S1378 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1951_ (
  .in1({ S1375, S257 }),
  .out1({ S1379 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1952_ (
  .in1({ S1378, S1376 }),
  .out1({ S1380 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1953_ (
  .in1({ S1379, S1377 }),
  .out1({ S1381 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1954_ (
  .in1({ S1267, new_datapath_addsubunit_in1_5 }),
  .out1({ S1382 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1955_ (
  .in1({ S1268, S5926 }),
  .out1({ S1383 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1956_ (
  .in1({ S1268, S1210 }),
  .out1({ S1384 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1957_ (
  .in1({ S1267, S1211 }),
  .out1({ S1385 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1958_ (
  .in1({ S1384, S1382 }),
  .out1({ S1386 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1959_ (
  .in1({ S1385, S1383 }),
  .out1({ S1387 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1960_ (
  .in1({ S1387, S265 }),
  .out1({ S1388 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1961_ (
  .in1({ S1386, S264 }),
  .out1({ S1389 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1962_ (
  .in1({ S1386, S264 }),
  .out1({ S1390 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1963_ (
  .in1({ S1387, S265 }),
  .out1({ S1391 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1964_ (
  .in1({ S1390, S1388 }),
  .out1({ S1392 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1965_ (
  .in1({ S1391, S1389 }),
  .out1({ S1393 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1966_ (
  .in1({ S1393, S1202 }),
  .out1({ S1394 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1967_ (
  .in1({ S1392, S1203 }),
  .out1({ S1395 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1968_ (
  .in1({ S1394, S1388 }),
  .out1({ S1396 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1969_ (
  .in1({ S1395, S1389 }),
  .out1({ S1397 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1970_ (
  .in1({ S1396, S1381 }),
  .out1({ S1398 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1971_ (
  .in1({ S1397, S1380 }),
  .out1({ S1399 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1972_ (
  .in1({ S1398, S1376 }),
  .out1({ S1400 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1973_ (
  .in1({ S1399, S1377 }),
  .out1({ S1401 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1974_ (
  .in1({ S1400, S1367 }),
  .out1({ S1402 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1975_ (
  .in1({ S1401, S1366 }),
  .out1({ S1403 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1976_ (
  .in1({ S1402, S1362 }),
  .out1({ S1404 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1977_ (
  .in1({ S1403, S1363 }),
  .out1({ S1405 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1978_ (
  .in1({ S1350, S240 }),
  .out1({ S1406 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1979_ (
  .in1({ S1351, S241 }),
  .out1({ S1407 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1980_ (
  .in1({ S1406, S1352 }),
  .out1({ S1408 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1981_ (
  .in1({ S1407, S1353 }),
  .out1({ S1409 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1982_ (
  .in1({ S1409, S1404 }),
  .out1({ S1410 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1983_ (
  .in1({ S1408, S1405 }),
  .out1({ S1411 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1984_ (
  .in1({ S1410, S1352 }),
  .out1({ S1412 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1985_ (
  .in1({ S1411, S1353 }),
  .out1({ S1413 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1986_ (
  .in1({ S1412, S1343 }),
  .out1({ S1414 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1987_ (
  .in1({ S1413, S1342 }),
  .out1({ S1415 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1988_ (
  .in1({ S1414, S1338 }),
  .out1({ S1416 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1989_ (
  .in1({ S1415, S1339 }),
  .out1({ S1417 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1990_ (
  .in1({ S1416, S1329 }),
  .out1({ S1418 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1991_ (
  .in1({ S1417, S1328 }),
  .out1({ S1419 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1992_ (
  .in1({ S1418, S1324 }),
  .out1({ S1420 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1993_ (
  .in1({ S1419, S1325 }),
  .out1({ S1421 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1994_ (
  .in1({ S1420, S1314 }),
  .out1({ S1422 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1995_ (
  .in1({ S1421, S1315 }),
  .out1({ S1423 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1996_ (
  .in1({ S1422, S1312 }),
  .out1({ S1424 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1997_ (
  .in1({ S1423, S1313 }),
  .out1({ S1425 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_1998_ (
  .in1({ S1424, S1302 }),
  .out1({ S1426 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_1999_ (
  .in1({ S1425, S1303 }),
  .out1({ S1427 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2000_ (
  .in1({ S1426, S1299 }),
  .out1({ S1428 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2001_ (
  .in1({ S1427, S1300 }),
  .out1({ S1429 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2002_ (
  .in1({ S1429, S1292 }),
  .out1({ S1430 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2003_ (
  .in1({ S1428, S1291 }),
  .out1({ S1431 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2004_ (
  .in1({ S1431, S1292 }),
  .out1({ S1432 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2005_ (
  .in1({ S1430, S1291 }),
  .out1({ S1433 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2006_ (
  .in1({ S1432, S1278 }),
  .out1({ S1434 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2007_ (
  .in1({ S1433, S1279 }),
  .out1({ S1435 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2008_ (
  .in1({ S1434, S1275 }),
  .out1({ S1436 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2009_ (
  .in1({ S1435, S1276 }),
  .out1({ S1437 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2010_ (
  .in1({ S214, new_datapath_multdivunit_1697_B_11 }),
  .out1({ S1438 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2011_ (
  .in1({ S1438, S1437 }),
  .out1({ S1439 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2012_ (
  .in1({ S1436, S217 }),
  .out1({ S1440 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2013_ (
  .in1({ S1440, S1439 }),
  .out1({ S1441 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2014_ (
  .in1({ S1441, S1259 }),
  .out1({ S1442 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2015_ (
  .in1({ S1442, new_datapath_multdivunit_1697_B_12 }),
  .out1({ S1443 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2016_ (
  .in1({ S1443 }),
  .out1({ S1444 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2017_ (
  .in1({ S1076, new_datapath_multdivunit_1697_B_11 }),
  .out1({ S1445 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2018_ (
  .in1({ S1445, S214 }),
  .out1({ S1446 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2019_ (
  .in1({ S1446 }),
  .out1({ S1447 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2020_ (
  .in1({ S1446, S1436 }),
  .out1({ S1448 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2021_ (
  .in1({ S1447, S1437 }),
  .out1({ S1449 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2022_ (
  .in1({ S1258, S217 }),
  .out1({ S1450 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2023_ (
  .in1({ S1259, S216 }),
  .out1({ S1451 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2024_ (
  .in1({ S1450, S1448 }),
  .out1({ S1452 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2025_ (
  .in1({ S1451, S1449 }),
  .out1({ S1453 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2026_ (
  .in1({ S1432, S1278 }),
  .out1({ S1454 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2027_ (
  .in1({ S1454, S1435 }),
  .out1({ S1455 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2028_ (
  .in1({ S1455, S1453 }),
  .out1({ S1456 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2029_ (
  .in1({ S1452, S1273 }),
  .out1({ S1457 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2030_ (
  .in1({ S1457, S1456 }),
  .out1({ S1458 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2031_ (
  .in1({ S1458 }),
  .out1({ S1459 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2032_ (
  .in1({ S1458, new_datapath_multdivunit_1697_B_11 }),
  .out1({ S1460 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2033_ (
  .in1({ S1459, S3445 }),
  .out1({ S1461 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2034_ (
  .in1({ S1458, new_datapath_multdivunit_1697_B_11 }),
  .out1({ S1462 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2035_ (
  .in1({ S1462, S1461 }),
  .out1({ S1463 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2036_ (
  .in1({ S1463 }),
  .out1({ S1464 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2037_ (
  .in1({ S1292, S1291 }),
  .out1({ S1465 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2038_ (
  .in1({ S1465, S1429 }),
  .out1({ S1466 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2039_ (
  .in1({ S1466 }),
  .out1({ S1467 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2040_ (
  .in1({ S1465, S1429 }),
  .out1({ S1468 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2041_ (
  .in1({ S1468, S1467 }),
  .out1({ S1469 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2042_ (
  .in1({ S1469, S1452 }),
  .out1({ S1470 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2043_ (
  .in1({ S1470 }),
  .out1({ S1471 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2044_ (
  .in1({ S1452, S1289 }),
  .out1({ S1472 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2045_ (
  .in1({ S1472 }),
  .out1({ S1473 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2046_ (
  .in1({ S1473, S1470 }),
  .out1({ S1474 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2047_ (
  .in1({ S1472, S1471 }),
  .out1({ S1475 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2048_ (
  .in1({ S1475, S3456 }),
  .out1({ S1476 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2049_ (
  .in1({ S1474, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S1477 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2050_ (
  .in1({ S1424, S1302 }),
  .out1({ S1478 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2051_ (
  .in1({ S1478, S1427 }),
  .out1({ S1479 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2052_ (
  .in1({ S1479, S1453 }),
  .out1({ S1480 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2053_ (
  .in1({ S1452, S1297 }),
  .out1({ S1481 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2054_ (
  .in1({ S1481, S1480 }),
  .out1({ S1482 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2055_ (
  .in1({ S1482 }),
  .out1({ S1483 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2056_ (
  .in1({ S1482, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S1484 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2057_ (
  .in1({ S1483, S3467 }),
  .out1({ S1485 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2058_ (
  .in1({ S1482, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S1486 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2059_ (
  .in1({ S1486, S1485 }),
  .out1({ S1487 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2060_ (
  .in1({ S1487 }),
  .out1({ S1488 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2061_ (
  .in1({ S1314, S1312 }),
  .out1({ S1489 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2062_ (
  .in1({ S1315, S1313 }),
  .out1({ S1490 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2063_ (
  .in1({ S1489, S1421 }),
  .out1({ S1491 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2064_ (
  .in1({ S1490, S1420 }),
  .out1({ S1492 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2065_ (
  .in1({ S1492, S1491 }),
  .out1({ S1493 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2066_ (
  .in1({ S1493, S1452 }),
  .out1({ S1494 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2067_ (
  .in1({ S1494 }),
  .out1({ S1495 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2068_ (
  .in1({ S1452, S1311 }),
  .out1({ S1496 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2069_ (
  .in1({ S1496 }),
  .out1({ S1497 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2070_ (
  .in1({ S1497, S1494 }),
  .out1({ S1498 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2071_ (
  .in1({ S1496, S1495 }),
  .out1({ S1499 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2072_ (
  .in1({ S1499, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S1500 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2073_ (
  .in1({ S1498, S3478 }),
  .out1({ S1501 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2074_ (
  .in1({ S1416, S1329 }),
  .out1({ S1502 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2075_ (
  .in1({ S1502, S1419 }),
  .out1({ S1503 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2076_ (
  .in1({ S1503, S1453 }),
  .out1({ S1504 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2077_ (
  .in1({ S1452, S1323 }),
  .out1({ S1505 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2078_ (
  .in1({ S1505, S1504 }),
  .out1({ S1506 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2079_ (
  .in1({ S1506 }),
  .out1({ S1507 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2080_ (
  .in1({ S1506, S229 }),
  .out1({ S1508 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2081_ (
  .in1({ S1507, S228 }),
  .out1({ S1509 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2082_ (
  .in1({ S1506, S229 }),
  .out1({ S1510 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2083_ (
  .in1({ S1510, S1509 }),
  .out1({ S1511 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2084_ (
  .in1({ S1511 }),
  .out1({ S1512 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2085_ (
  .in1({ S1413, S1342 }),
  .out1({ S1513 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2086_ (
  .in1({ S1513, S1414 }),
  .out1({ S1514 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2087_ (
  .in1({ S1514, S1452 }),
  .out1({ S1515 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2088_ (
  .in1({ S1515 }),
  .out1({ S1516 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2089_ (
  .in1({ S1452, S1337 }),
  .out1({ S1517 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2090_ (
  .in1({ S1517 }),
  .out1({ S1518 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2091_ (
  .in1({ S1518, S1515 }),
  .out1({ S1519 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2092_ (
  .in1({ S1517, S1516 }),
  .out1({ S1520 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2093_ (
  .in1({ S1519, S202 }),
  .out1({ S1521 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2094_ (
  .in1({ S1520, S203 }),
  .out1({ S1522 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2095_ (
  .in1({ S1408, S1405 }),
  .out1({ S1523 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2096_ (
  .in1({ S1523, S1410 }),
  .out1({ S1524 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2097_ (
  .in1({ S1524, S1452 }),
  .out1({ S1525 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2098_ (
  .in1({ S1453, S1350 }),
  .out1({ S1526 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2099_ (
  .in1({ S1526, S1525 }),
  .out1({ S1527 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2100_ (
  .in1({ S1527 }),
  .out1({ S1528 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2101_ (
  .in1({ S1528, S209 }),
  .out1({ S1529 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2102_ (
  .in1({ S1527, S208 }),
  .out1({ S1530 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2103_ (
  .in1({ S1453, S1360 }),
  .out1({ S1531 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2104_ (
  .in1({ S1452, S1361 }),
  .out1({ S1532 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2105_ (
  .in1({ S1401, S1366 }),
  .out1({ S1533 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2106_ (
  .in1({ S1533, S1402 }),
  .out1({ S1534 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2107_ (
  .in1({ S1534, S1452 }),
  .out1({ S1535 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2108_ (
  .in1({ S1535 }),
  .out1({ S1536 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2109_ (
  .in1({ S1535, S1531 }),
  .out1({ S1537 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2110_ (
  .in1({ S1536, S1532 }),
  .out1({ S1538 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2111_ (
  .in1({ S1538, S241 }),
  .out1({ S1539 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2112_ (
  .in1({ S1537, S240 }),
  .out1({ S1540 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2113_ (
  .in1({ S1537, S240 }),
  .out1({ S1541 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2114_ (
  .in1({ S1538, S241 }),
  .out1({ S1542 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2115_ (
  .in1({ S1541, S1539 }),
  .out1({ S1543 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2116_ (
  .in1({ S1542, S1540 }),
  .out1({ S1544 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2117_ (
  .in1({ S1396, S1381 }),
  .out1({ S1545 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2118_ (
  .in1({ S1545, S1399 }),
  .out1({ S1546 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2119_ (
  .in1({ S1546, S1453 }),
  .out1({ S1547 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2120_ (
  .in1({ S1452, S1375 }),
  .out1({ S1548 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2121_ (
  .in1({ S1548, S1547 }),
  .out1({ S1549 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2122_ (
  .in1({ S1549 }),
  .out1({ S1550 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2123_ (
  .in1({ S1549, S249 }),
  .out1({ S1551 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2124_ (
  .in1({ S1550, S248 }),
  .out1({ S1552 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2125_ (
  .in1({ S1549, S249 }),
  .out1({ S1553 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2126_ (
  .in1({ S1553, S1552 }),
  .out1({ S1554 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2127_ (
  .in1({ S1554 }),
  .out1({ S1555 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2128_ (
  .in1({ S1392, S1203 }),
  .out1({ S1556 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2129_ (
  .in1({ S1556, S1394 }),
  .out1({ S1557 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2130_ (
  .in1({ S1557, S1452 }),
  .out1({ S1558 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2131_ (
  .in1({ S1453, S1386 }),
  .out1({ S1559 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2132_ (
  .in1({ S1559, S1558 }),
  .out1({ S1560 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2133_ (
  .in1({ S1560 }),
  .out1({ S1561 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2134_ (
  .in1({ S1561, S257 }),
  .out1({ S1562 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2135_ (
  .in1({ S1560, S256 }),
  .out1({ S1563 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2136_ (
  .in1({ S1560, S256 }),
  .out1({ S1564 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2137_ (
  .in1({ S1561, S257 }),
  .out1({ S1565 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2138_ (
  .in1({ S1452, S270 }),
  .out1({ S1566 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2139_ (
  .in1({ S1453, S271 }),
  .out1({ S1567 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2140_ (
  .in1({ S1566, S5936 }),
  .out1({ S1568 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2141_ (
  .in1({ S1567, new_datapath_addsubunit_in1_4 }),
  .out1({ S1569 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2142_ (
  .in1({ S1452, S1203 }),
  .out1({ S1570 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2143_ (
  .in1({ S1453, S1202 }),
  .out1({ S1571 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2144_ (
  .in1({ S1570, S1568 }),
  .out1({ S1572 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2145_ (
  .in1({ S1571, S1569 }),
  .out1({ S1573 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2146_ (
  .in1({ S1572, S265 }),
  .out1({ S1574 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2147_ (
  .in1({ S1573, S264 }),
  .out1({ S1575 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2148_ (
  .in1({ S1573, S264 }),
  .out1({ S1576 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2149_ (
  .in1({ S1572, S265 }),
  .out1({ S1577 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2150_ (
  .in1({ S1576, S1574 }),
  .out1({ S1578 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2151_ (
  .in1({ S1577, S1575 }),
  .out1({ S1579 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2152_ (
  .in1({ S270, new_datapath_addsubunit_in1_3 }),
  .out1({ S1580 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2153_ (
  .in1({ S271, S5947 }),
  .out1({ S1581 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2154_ (
  .in1({ S1580, S1579 }),
  .out1({ S1582 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2155_ (
  .in1({ S1581, S1578 }),
  .out1({ S1583 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2156_ (
  .in1({ S1582, S1574 }),
  .out1({ S1584 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2157_ (
  .in1({ S1583, S1575 }),
  .out1({ S1585 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2158_ (
  .in1({ S1584, S1564 }),
  .out1({ S1586 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2159_ (
  .in1({ S1585, S1565 }),
  .out1({ S1587 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2160_ (
  .in1({ S1586, S1562 }),
  .out1({ S1588 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2161_ (
  .in1({ S1587, S1563 }),
  .out1({ S1589 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2162_ (
  .in1({ S1588, S1554 }),
  .out1({ S1590 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2163_ (
  .in1({ S1589, S1555 }),
  .out1({ S1591 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2164_ (
  .in1({ S1590, S1551 }),
  .out1({ S1592 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2165_ (
  .in1({ S1591, S1552 }),
  .out1({ S1593 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2166_ (
  .in1({ S1592, S1544 }),
  .out1({ S1594 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2167_ (
  .in1({ S1593, S1543 }),
  .out1({ S1595 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2168_ (
  .in1({ S1594, S1539 }),
  .out1({ S1596 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2169_ (
  .in1({ S1595, S1540 }),
  .out1({ S1597 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2170_ (
  .in1({ S1527, S208 }),
  .out1({ S1598 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2171_ (
  .in1({ S1598, S1529 }),
  .out1({ S1599 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2172_ (
  .in1({ S1599 }),
  .out1({ S1600 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2173_ (
  .in1({ S1600, S1596 }),
  .out1({ S1601 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2174_ (
  .in1({ S1599, S1597 }),
  .out1({ S1602 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2175_ (
  .in1({ S1601, S1529 }),
  .out1({ S1603 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2176_ (
  .in1({ S1602, S1530 }),
  .out1({ S1604 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2177_ (
  .in1({ S1604, S1522 }),
  .out1({ S1605 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2178_ (
  .in1({ S1603, S1521 }),
  .out1({ S1606 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2179_ (
  .in1({ S1606, S1522 }),
  .out1({ S1607 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2180_ (
  .in1({ S1605, S1521 }),
  .out1({ S1608 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2181_ (
  .in1({ S1607, S1511 }),
  .out1({ S1609 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2182_ (
  .in1({ S1608, S1512 }),
  .out1({ S1610 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2183_ (
  .in1({ S1609, S1508 }),
  .out1({ S1611 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2184_ (
  .in1({ S1610, S1509 }),
  .out1({ S1612 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2185_ (
  .in1({ S1611, S1501 }),
  .out1({ S1613 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2186_ (
  .in1({ S1612, S1500 }),
  .out1({ S1614 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2187_ (
  .in1({ S1613, S1500 }),
  .out1({ S1615 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2188_ (
  .in1({ S1614, S1501 }),
  .out1({ S1616 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2189_ (
  .in1({ S1615, S1487 }),
  .out1({ S1617 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2190_ (
  .in1({ S1616, S1488 }),
  .out1({ S1618 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2191_ (
  .in1({ S1617, S1484 }),
  .out1({ S1619 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2192_ (
  .in1({ S1618, S1485 }),
  .out1({ S1620 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2193_ (
  .in1({ S1620, S1477 }),
  .out1({ S1621 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2194_ (
  .in1({ S1619, S1476 }),
  .out1({ S1622 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2195_ (
  .in1({ S1621, S1476 }),
  .out1({ S1623 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2196_ (
  .in1({ S1622, S1477 }),
  .out1({ S1624 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2197_ (
  .in1({ S1624, S1463 }),
  .out1({ S1625 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2198_ (
  .in1({ S1623, S1464 }),
  .out1({ S1626 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2199_ (
  .in1({ S1625, S1460 }),
  .out1({ S1627 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2200_ (
  .in1({ S1626, S1461 }),
  .out1({ S1628 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2201_ (
  .in1({ S1628, S1443 }),
  .out1({ S1629 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2202_ (
  .in1({ S1627, S1444 }),
  .out1({ S1630 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2203_ (
  .in1({ S1258, new_datapath_multdivunit_1697_B_12 }),
  .out1({ S1631 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2204_ (
  .in1({ S1631, S212 }),
  .out1({ S1632 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2205_ (
  .in1({ S1632 }),
  .out1({ S1633 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2206_ (
  .in1({ S1632, S1629 }),
  .out1({ S1634 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2207_ (
  .in1({ S1633, S1630 }),
  .out1({ S1635 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2208_ (
  .in1({ S1624, S1463 }),
  .out1({ S1636 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2209_ (
  .in1({ S1636, S1626 }),
  .out1({ S1637 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2210_ (
  .in1({ S1637, S1634 }),
  .out1({ S1638 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2211_ (
  .in1({ S1635, S1458 }),
  .out1({ S1639 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2212_ (
  .in1({ S1639, S1638 }),
  .out1({ S1640 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2213_ (
  .in1({ S1640 }),
  .out1({ S1641 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2214_ (
  .in1({ S1640, new_datapath_multdivunit_1697_B_12 }),
  .out1({ S1642 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2215_ (
  .in1({ S1641, S3434 }),
  .out1({ S1643 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2216_ (
  .in1({ S1640, new_datapath_multdivunit_1697_B_12 }),
  .out1({ S1644 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2217_ (
  .in1({ S1644, S1643 }),
  .out1({ S1645 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2218_ (
  .in1({ S1645 }),
  .out1({ S1646 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2219_ (
  .in1({ S1477, S1476 }),
  .out1({ S1647 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2220_ (
  .in1({ S1647, S1620 }),
  .out1({ S1648 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2221_ (
  .in1({ S1648 }),
  .out1({ S1649 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2222_ (
  .in1({ S1647, S1620 }),
  .out1({ S1650 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2223_ (
  .in1({ S1650 }),
  .out1({ S1651 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2224_ (
  .in1({ S1651, S1648 }),
  .out1({ S1652 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2225_ (
  .in1({ S1650, S1649 }),
  .out1({ S1653 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2226_ (
  .in1({ S1652, S1635 }),
  .out1({ S1654 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2227_ (
  .in1({ S1653, S1634 }),
  .out1({ S1655 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2228_ (
  .in1({ S1634, S1475 }),
  .out1({ S1656 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2229_ (
  .in1({ S1635, S1474 }),
  .out1({ S1657 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2230_ (
  .in1({ S1656, S1654 }),
  .out1({ S1658 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2231_ (
  .in1({ S1657, S1655 }),
  .out1({ S1659 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2232_ (
  .in1({ S1659, new_datapath_multdivunit_1697_B_11 }),
  .out1({ S1660 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2233_ (
  .in1({ S1658, S3445 }),
  .out1({ S1661 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2234_ (
  .in1({ S1658, S3445 }),
  .out1({ S1662 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2235_ (
  .in1({ S1659, new_datapath_multdivunit_1697_B_11 }),
  .out1({ S1663 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2236_ (
  .in1({ S1615, S1487 }),
  .out1({ S1664 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2237_ (
  .in1({ S1664, S1618 }),
  .out1({ S1665 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2238_ (
  .in1({ S1665, S1634 }),
  .out1({ S1666 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2239_ (
  .in1({ S1635, S1482 }),
  .out1({ S1667 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2240_ (
  .in1({ S1667, S1666 }),
  .out1({ S1668 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2241_ (
  .in1({ S1668 }),
  .out1({ S1669 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2242_ (
  .in1({ S1668, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S1670 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2243_ (
  .in1({ S1669, S3456 }),
  .out1({ S1671 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2244_ (
  .in1({ S1668, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S1672 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2245_ (
  .in1({ S1672 }),
  .out1({ S1673 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2246_ (
  .in1({ S1673, S1670 }),
  .out1({ S1674 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2247_ (
  .in1({ S1672, S1671 }),
  .out1({ S1675 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2248_ (
  .in1({ S1501, S1500 }),
  .out1({ S1676 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2249_ (
  .in1({ S1676, S1612 }),
  .out1({ S1677 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2250_ (
  .in1({ S1677 }),
  .out1({ S1678 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2251_ (
  .in1({ S1676, S1612 }),
  .out1({ S1679 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2252_ (
  .in1({ S1679 }),
  .out1({ S1680 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2253_ (
  .in1({ S1680, S1677 }),
  .out1({ S1681 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2254_ (
  .in1({ S1679, S1678 }),
  .out1({ S1682 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2255_ (
  .in1({ S1681, S1635 }),
  .out1({ S1683 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2256_ (
  .in1({ S1682, S1634 }),
  .out1({ S1684 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2257_ (
  .in1({ S1634, S1498 }),
  .out1({ S1685 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2258_ (
  .in1({ S1635, S1499 }),
  .out1({ S1686 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2259_ (
  .in1({ S1685, S1683 }),
  .out1({ S1687 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2260_ (
  .in1({ S1686, S1684 }),
  .out1({ S1688 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2261_ (
  .in1({ S1687, S3467 }),
  .out1({ S1689 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2262_ (
  .in1({ S1688, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S1690 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2263_ (
  .in1({ S1607, S1511 }),
  .out1({ S1691 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2264_ (
  .in1({ S1691, S1610 }),
  .out1({ S1692 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2265_ (
  .in1({ S1692, S1634 }),
  .out1({ S1693 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2266_ (
  .in1({ S1635, S1506 }),
  .out1({ S1694 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2267_ (
  .in1({ S1694, S1693 }),
  .out1({ S1695 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2268_ (
  .in1({ S1695 }),
  .out1({ S1696 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2269_ (
  .in1({ S1695, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S1697 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2270_ (
  .in1({ S1696, S3478 }),
  .out1({ S1698 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2271_ (
  .in1({ S1695, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S1699 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2272_ (
  .in1({ S1699, S1698 }),
  .out1({ S1700 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2273_ (
  .in1({ S1700 }),
  .out1({ S1701 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2274_ (
  .in1({ S1522, S1521 }),
  .out1({ S1702 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2275_ (
  .in1({ S1702, S1603 }),
  .out1({ S1703 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2276_ (
  .in1({ S1703 }),
  .out1({ S1704 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2277_ (
  .in1({ S1702, S1603 }),
  .out1({ S1705 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2278_ (
  .in1({ S1705, S1704 }),
  .out1({ S1706 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2279_ (
  .in1({ S1706, S1635 }),
  .out1({ S1707 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2280_ (
  .in1({ S1634, S1519 }),
  .out1({ S1708 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2281_ (
  .in1({ S1708, S1707 }),
  .out1({ S1709 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2282_ (
  .in1({ S1709 }),
  .out1({ S1710 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2283_ (
  .in1({ S1709, S228 }),
  .out1({ S1711 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2284_ (
  .in1({ S1710, S229 }),
  .out1({ S1712 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2285_ (
  .in1({ S1599, S1597 }),
  .out1({ S1713 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2286_ (
  .in1({ S1713, S1601 }),
  .out1({ S1714 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2287_ (
  .in1({ S1714, S1635 }),
  .out1({ S1715 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2288_ (
  .in1({ S1634, S1527 }),
  .out1({ S1716 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2289_ (
  .in1({ S1716, S1715 }),
  .out1({ S1717 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2290_ (
  .in1({ S1717 }),
  .out1({ S1718 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2291_ (
  .in1({ S1718, S203 }),
  .out1({ S1719 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2292_ (
  .in1({ S1719 }),
  .out1({ S1720 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2293_ (
  .in1({ S1593, S1543 }),
  .out1({ S1721 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2294_ (
  .in1({ S1721 }),
  .out1({ S1722 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2295_ (
  .in1({ S1721, S1594 }),
  .out1({ S1723 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2296_ (
  .in1({ S1722, S1595 }),
  .out1({ S1724 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2297_ (
  .in1({ S1723, S1635 }),
  .out1({ S1725 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2298_ (
  .in1({ S1724, S1634 }),
  .out1({ S1726 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2299_ (
  .in1({ S1634, S1537 }),
  .out1({ S1727 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2300_ (
  .in1({ S1635, S1538 }),
  .out1({ S1728 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2301_ (
  .in1({ S1727, S1725 }),
  .out1({ S1729 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2302_ (
  .in1({ S1728, S1726 }),
  .out1({ S1730 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2303_ (
  .in1({ S1730, S209 }),
  .out1({ S1731 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2304_ (
  .in1({ S1729, S208 }),
  .out1({ S1732 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2305_ (
  .in1({ S1729, S208 }),
  .out1({ S1733 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2306_ (
  .in1({ S1733, S1731 }),
  .out1({ S1734 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2307_ (
  .in1({ S1734 }),
  .out1({ S1735 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2308_ (
  .in1({ S1588, S1554 }),
  .out1({ S1736 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2309_ (
  .in1({ S1736, S1591 }),
  .out1({ S1737 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2310_ (
  .in1({ S1737, S1634 }),
  .out1({ S1738 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2311_ (
  .in1({ S1635, S1549 }),
  .out1({ S1739 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2312_ (
  .in1({ S1739, S1738 }),
  .out1({ S1740 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2313_ (
  .in1({ S1740 }),
  .out1({ S1741 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2314_ (
  .in1({ S1741, S240 }),
  .out1({ S1742 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2315_ (
  .in1({ S1742 }),
  .out1({ S1743 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2316_ (
  .in1({ S1740, S241 }),
  .out1({ S1744 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2317_ (
  .in1({ S1744, S1742 }),
  .out1({ S1745 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2318_ (
  .in1({ S1745 }),
  .out1({ S1746 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2319_ (
  .in1({ S1564, S1562 }),
  .out1({ S1747 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2320_ (
  .in1({ S1565, S1563 }),
  .out1({ S1748 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2321_ (
  .in1({ S1747, S1584 }),
  .out1({ S1749 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2322_ (
  .in1({ S1748, S1585 }),
  .out1({ S1750 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2323_ (
  .in1({ S1750, S1749 }),
  .out1({ S1751 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2324_ (
  .in1({ S1751, S1634 }),
  .out1({ S1752 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2325_ (
  .in1({ S1635, S1560 }),
  .out1({ S1753 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2326_ (
  .in1({ S1753, S1752 }),
  .out1({ S1754 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2327_ (
  .in1({ S1754 }),
  .out1({ S1755 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2328_ (
  .in1({ S1755, S249 }),
  .out1({ S1756 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2329_ (
  .in1({ S1756 }),
  .out1({ S1757 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2330_ (
  .in1({ S1754, S248 }),
  .out1({ S1758 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2331_ (
  .in1({ S1758, S1756 }),
  .out1({ S1759 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2332_ (
  .in1({ S1759 }),
  .out1({ S1760 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2333_ (
  .in1({ S1581, S1578 }),
  .out1({ S1761 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2334_ (
  .in1({ S1580, S1579 }),
  .out1({ S1762 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2335_ (
  .in1({ S1761, S1582 }),
  .out1({ S1763 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2336_ (
  .in1({ S1762, S1583 }),
  .out1({ S1764 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2337_ (
  .in1({ S1763, S1635 }),
  .out1({ S1765 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2338_ (
  .in1({ S1764, S1634 }),
  .out1({ S1766 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2339_ (
  .in1({ S1634, S1573 }),
  .out1({ S1767 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2340_ (
  .in1({ S1635, S1572 }),
  .out1({ S1768 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2341_ (
  .in1({ S1767, S1765 }),
  .out1({ S1769 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2342_ (
  .in1({ S1768, S1766 }),
  .out1({ S1770 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2343_ (
  .in1({ S1770, S257 }),
  .out1({ S1771 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2344_ (
  .in1({ S1769, S256 }),
  .out1({ S1772 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2345_ (
  .in1({ S1769, S256 }),
  .out1({ S1773 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2346_ (
  .in1({ S1770, S257 }),
  .out1({ S1774 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2347_ (
  .in1({ S1773, S1771 }),
  .out1({ S1775 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2348_ (
  .in1({ S1774, S1772 }),
  .out1({ S1776 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2349_ (
  .in1({ S1635, S270 }),
  .out1({ S1777 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2350_ (
  .in1({ S1634, S271 }),
  .out1({ S1778 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2351_ (
  .in1({ S1777, S5947 }),
  .out1({ S1779 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2352_ (
  .in1({ S1778, new_datapath_addsubunit_in1_3 }),
  .out1({ S1780 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2353_ (
  .in1({ S1635, S1581 }),
  .out1({ S1781 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2354_ (
  .in1({ S1634, S1580 }),
  .out1({ S1782 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2355_ (
  .in1({ S1781, S1779 }),
  .out1({ S1783 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2356_ (
  .in1({ S1782, S1780 }),
  .out1({ S1784 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2357_ (
  .in1({ S1783, S265 }),
  .out1({ S1785 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2358_ (
  .in1({ S1784, S264 }),
  .out1({ S1786 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2359_ (
  .in1({ S270, new_datapath_addsubunit_in1_2 }),
  .out1({ S1787 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2360_ (
  .in1({ S271, S5957 }),
  .out1({ S1788 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2361_ (
  .in1({ S1784, S264 }),
  .out1({ S1789 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2362_ (
  .in1({ S1783, S265 }),
  .out1({ S1790 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2363_ (
  .in1({ S1789, S1785 }),
  .out1({ S1791 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2364_ (
  .in1({ S1790, S1786 }),
  .out1({ S1792 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2365_ (
  .in1({ S1792, S1787 }),
  .out1({ S1793 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2366_ (
  .in1({ S1791, S1788 }),
  .out1({ S1794 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2367_ (
  .in1({ S1793, S1785 }),
  .out1({ S1795 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2368_ (
  .in1({ S1794, S1786 }),
  .out1({ S1796 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2369_ (
  .in1({ S1795, S1776 }),
  .out1({ S1797 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2370_ (
  .in1({ S1796, S1775 }),
  .out1({ S1798 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2371_ (
  .in1({ S1797, S1771 }),
  .out1({ S1799 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2372_ (
  .in1({ S1798, S1772 }),
  .out1({ S1800 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2373_ (
  .in1({ S1799, S1760 }),
  .out1({ S1801 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2374_ (
  .in1({ S1800, S1759 }),
  .out1({ S1802 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2375_ (
  .in1({ S1801, S1756 }),
  .out1({ S1803 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2376_ (
  .in1({ S1802, S1757 }),
  .out1({ S1804 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2377_ (
  .in1({ S1803, S1745 }),
  .out1({ S1805 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2378_ (
  .in1({ S1804, S1746 }),
  .out1({ S1806 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2379_ (
  .in1({ S1805, S1743 }),
  .out1({ S1807 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2380_ (
  .in1({ S1806, S1742 }),
  .out1({ S1808 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2381_ (
  .in1({ S1807, S1735 }),
  .out1({ S1809 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2382_ (
  .in1({ S1808, S1734 }),
  .out1({ S1810 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2383_ (
  .in1({ S1809, S1731 }),
  .out1({ S1811 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2384_ (
  .in1({ S1810, S1732 }),
  .out1({ S1812 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2385_ (
  .in1({ S1717, S202 }),
  .out1({ S1813 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2386_ (
  .in1({ S1813, S1719 }),
  .out1({ S1814 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2387_ (
  .in1({ S1814 }),
  .out1({ S1815 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2388_ (
  .in1({ S1815, S1811 }),
  .out1({ S1816 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2389_ (
  .in1({ S1814, S1812 }),
  .out1({ S1817 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2390_ (
  .in1({ S1816, S1719 }),
  .out1({ S1818 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2391_ (
  .in1({ S1817, S1720 }),
  .out1({ S1819 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2392_ (
  .in1({ S1819, S1712 }),
  .out1({ S1820 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2393_ (
  .in1({ S1818, S1711 }),
  .out1({ S1821 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2394_ (
  .in1({ S1821, S1712 }),
  .out1({ S1822 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2395_ (
  .in1({ S1820, S1711 }),
  .out1({ S1823 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2396_ (
  .in1({ S1822, S1700 }),
  .out1({ S1824 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2397_ (
  .in1({ S1823, S1701 }),
  .out1({ S1825 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2398_ (
  .in1({ S1824, S1697 }),
  .out1({ S1826 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2399_ (
  .in1({ S1825, S1698 }),
  .out1({ S1827 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2400_ (
  .in1({ S1827, S1690 }),
  .out1({ S1828 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2401_ (
  .in1({ S1826, S1689 }),
  .out1({ S1829 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2402_ (
  .in1({ S1829, S1690 }),
  .out1({ S1830 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2403_ (
  .in1({ S1828, S1689 }),
  .out1({ S1831 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2404_ (
  .in1({ S1830, S1675 }),
  .out1({ S1832 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2405_ (
  .in1({ S1831, S1674 }),
  .out1({ S1833 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2406_ (
  .in1({ S1832, S1670 }),
  .out1({ S1834 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2407_ (
  .in1({ S1833, S1671 }),
  .out1({ S1835 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2408_ (
  .in1({ S1834, S1662 }),
  .out1({ S1836 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2409_ (
  .in1({ S1835, S1663 }),
  .out1({ S1837 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2410_ (
  .in1({ S1836, S1660 }),
  .out1({ S1838 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2411_ (
  .in1({ S1837, S1661 }),
  .out1({ S1839 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2412_ (
  .in1({ S1838, S1645 }),
  .out1({ S1840 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2413_ (
  .in1({ S1839, S1646 }),
  .out1({ S1841 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2414_ (
  .in1({ S1840, S1642 }),
  .out1({ S1842 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2415_ (
  .in1({ S1841, S1643 }),
  .out1({ S1843 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2416_ (
  .in1({ S212, new_datapath_multdivunit_1697_B_12 }),
  .out1({ S1844 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2417_ (
  .in1({ S1627, S214 }),
  .out1({ S1845 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2418_ (
  .in1({ S1844, S1627 }),
  .out1({ S1846 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2419_ (
  .in1({ S1846, S1442 }),
  .out1({ S1847 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2420_ (
  .in1({ S1847, S1845 }),
  .out1({ S1848 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2421_ (
  .in1({ S1848, new_datapath_multdivunit_1697_B_13 }),
  .out1({ S1849 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2422_ (
  .in1({ S1849 }),
  .out1({ S1850 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2423_ (
  .in1({ S1849, S1843 }),
  .out1({ S1851 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2424_ (
  .in1({ S1850, S1842 }),
  .out1({ S1852 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2425_ (
  .in1({ S1442, new_datapath_multdivunit_1697_B_13 }),
  .out1({ S1853 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2426_ (
  .in1({ S1853, S210 }),
  .out1({ S1854 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2427_ (
  .in1({ S1854 }),
  .out1({ S1855 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2428_ (
  .in1({ S1854, S1851 }),
  .out1({ S1856 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2429_ (
  .in1({ S1855, S1852 }),
  .out1({ S1857 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2430_ (
  .in1({ S1838, S1645 }),
  .out1({ S1858 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2431_ (
  .in1({ S1858, S1841 }),
  .out1({ S1859 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2432_ (
  .in1({ S1859, S1856 }),
  .out1({ S1860 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2433_ (
  .in1({ S1857, S1640 }),
  .out1({ S1861 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2434_ (
  .in1({ S1861, S1860 }),
  .out1({ S1862 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2435_ (
  .in1({ S1862 }),
  .out1({ S1863 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2436_ (
  .in1({ S1862, new_datapath_multdivunit_1697_B_13 }),
  .out1({ S1864 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2437_ (
  .in1({ S1863, S3423 }),
  .out1({ S1865 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2438_ (
  .in1({ S1862, new_datapath_multdivunit_1697_B_13 }),
  .out1({ S1866 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2439_ (
  .in1({ S1866, S1865 }),
  .out1({ S1867 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2440_ (
  .in1({ S1867 }),
  .out1({ S1868 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2441_ (
  .in1({ S1662, S1660 }),
  .out1({ S1869 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2442_ (
  .in1({ S1663, S1661 }),
  .out1({ S1870 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2443_ (
  .in1({ S1869, S1835 }),
  .out1({ S1871 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2444_ (
  .in1({ S1870, S1834 }),
  .out1({ S1872 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2445_ (
  .in1({ S1872, S1871 }),
  .out1({ S1873 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2446_ (
  .in1({ S1873, S1857 }),
  .out1({ S1874 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2447_ (
  .in1({ S1874 }),
  .out1({ S1875 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2448_ (
  .in1({ S1857, S1659 }),
  .out1({ S1876 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2449_ (
  .in1({ S1876 }),
  .out1({ S1877 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2450_ (
  .in1({ S1877, S1874 }),
  .out1({ S1878 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2451_ (
  .in1({ S1876, S1875 }),
  .out1({ S1879 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2452_ (
  .in1({ S1878, S3434 }),
  .out1({ S1880 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2453_ (
  .in1({ S1879, new_datapath_multdivunit_1697_B_12 }),
  .out1({ S1881 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2454_ (
  .in1({ S1830, S1675 }),
  .out1({ S1882 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2455_ (
  .in1({ S1882 }),
  .out1({ S1883 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2456_ (
  .in1({ S1883, S1832 }),
  .out1({ S1884 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2457_ (
  .in1({ S1884, S1857 }),
  .out1({ S1885 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2458_ (
  .in1({ S1885 }),
  .out1({ S1886 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2459_ (
  .in1({ S1857, S1668 }),
  .out1({ S1887 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2460_ (
  .in1({ S1887 }),
  .out1({ S1888 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2461_ (
  .in1({ S1888, S1885 }),
  .out1({ S1889 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2462_ (
  .in1({ S1887, S1886 }),
  .out1({ S1890 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2463_ (
  .in1({ S1890, new_datapath_multdivunit_1697_B_11 }),
  .out1({ S1891 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2464_ (
  .in1({ S1891 }),
  .out1({ S1892 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2465_ (
  .in1({ S1890, new_datapath_multdivunit_1697_B_11 }),
  .out1({ S1893 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2466_ (
  .in1({ S1893 }),
  .out1({ S1894 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2467_ (
  .in1({ S1894, S1891 }),
  .out1({ S1895 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2468_ (
  .in1({ S1895 }),
  .out1({ S1896 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2469_ (
  .in1({ S1690, S1689 }),
  .out1({ S1897 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2470_ (
  .in1({ S1897, S1826 }),
  .out1({ S1898 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2471_ (
  .in1({ S1898 }),
  .out1({ S1899 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2472_ (
  .in1({ S1897, S1826 }),
  .out1({ S1900 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2473_ (
  .in1({ S1900, S1899 }),
  .out1({ S1901 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2474_ (
  .in1({ S1901, S1857 }),
  .out1({ S1902 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2475_ (
  .in1({ S1902 }),
  .out1({ S1903 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2476_ (
  .in1({ S1857, S1688 }),
  .out1({ S1904 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2477_ (
  .in1({ S1904 }),
  .out1({ S1905 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2478_ (
  .in1({ S1905, S1902 }),
  .out1({ S1906 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2479_ (
  .in1({ S1904, S1903 }),
  .out1({ S1907 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2480_ (
  .in1({ S1906, S3456 }),
  .out1({ S1908 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2481_ (
  .in1({ S1907, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S1909 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2482_ (
  .in1({ S1822, S1700 }),
  .out1({ S1910 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2483_ (
  .in1({ S1910, S1825 }),
  .out1({ S1911 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2484_ (
  .in1({ S1911, S1856 }),
  .out1({ S1912 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2485_ (
  .in1({ S1857, S1695 }),
  .out1({ S1913 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2486_ (
  .in1({ S1913, S1912 }),
  .out1({ S1914 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2487_ (
  .in1({ S1914 }),
  .out1({ S1915 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2488_ (
  .in1({ S1914, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S1916 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2489_ (
  .in1({ S1915, S3467 }),
  .out1({ S1917 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2490_ (
  .in1({ S1914, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S1918 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2491_ (
  .in1({ S1918, S1917 }),
  .out1({ S1919 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2492_ (
  .in1({ S1919 }),
  .out1({ S1920 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2493_ (
  .in1({ S1712, S1711 }),
  .out1({ S1921 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2494_ (
  .in1({ S1921, S1818 }),
  .out1({ S1922 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2495_ (
  .in1({ S1922 }),
  .out1({ S1923 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2496_ (
  .in1({ S1921, S1818 }),
  .out1({ S1924 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2497_ (
  .in1({ S1924, S1923 }),
  .out1({ S1925 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2498_ (
  .in1({ S1925, S1857 }),
  .out1({ S1926 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2499_ (
  .in1({ S1857, S1710 }),
  .out1({ S1927 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2500_ (
  .in1({ S1927 }),
  .out1({ S1928 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2501_ (
  .in1({ S1928, S1926 }),
  .out1({ S1929 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2502_ (
  .in1({ S1929 }),
  .out1({ S1930 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2503_ (
  .in1({ S1929, S3478 }),
  .out1({ S1931 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2504_ (
  .in1({ S1930, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S1932 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2505_ (
  .in1({ S1814, S1812 }),
  .out1({ S1933 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2506_ (
  .in1({ S1933, S1816 }),
  .out1({ S1934 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2507_ (
  .in1({ S1934, S1857 }),
  .out1({ S1935 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2508_ (
  .in1({ S1856, S1717 }),
  .out1({ S1936 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2509_ (
  .in1({ S1936, S1935 }),
  .out1({ S1937 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2510_ (
  .in1({ S1937 }),
  .out1({ S1938 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2511_ (
  .in1({ S1938, S229 }),
  .out1({ S1939 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2512_ (
  .in1({ S1939 }),
  .out1({ S1940 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2513_ (
  .in1({ S1937, S228 }),
  .out1({ S1941 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2514_ (
  .in1({ S1941, S1939 }),
  .out1({ S1942 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2515_ (
  .in1({ S1942 }),
  .out1({ S1943 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2516_ (
  .in1({ S1857, S1730 }),
  .out1({ S1944 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2517_ (
  .in1({ S1944 }),
  .out1({ S1945 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2518_ (
  .in1({ S1808, S1734 }),
  .out1({ S1946 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2519_ (
  .in1({ S1946, S1809 }),
  .out1({ S1947 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2520_ (
  .in1({ S1947, S1857 }),
  .out1({ S1948 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2521_ (
  .in1({ S1948 }),
  .out1({ S1949 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2522_ (
  .in1({ S1948, S1945 }),
  .out1({ S1950 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2523_ (
  .in1({ S1949, S1944 }),
  .out1({ S1951 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2524_ (
  .in1({ S1951, S203 }),
  .out1({ S1952 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2525_ (
  .in1({ S1950, S202 }),
  .out1({ S1953 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2526_ (
  .in1({ S1803, S1745 }),
  .out1({ S1954 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2527_ (
  .in1({ S1954, S1806 }),
  .out1({ S1955 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2528_ (
  .in1({ S1955, S1856 }),
  .out1({ S1956 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2529_ (
  .in1({ S1857, S1740 }),
  .out1({ S1957 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2530_ (
  .in1({ S1957, S1956 }),
  .out1({ S1958 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2531_ (
  .in1({ S1958 }),
  .out1({ S1959 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2532_ (
  .in1({ S1959, S208 }),
  .out1({ S1960 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2533_ (
  .in1({ S1960 }),
  .out1({ S1961 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2534_ (
  .in1({ S1958, S209 }),
  .out1({ S1962 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2535_ (
  .in1({ S1962, S1960 }),
  .out1({ S1963 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2536_ (
  .in1({ S1963 }),
  .out1({ S1964 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2537_ (
  .in1({ S1800, S1759 }),
  .out1({ S1965 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2538_ (
  .in1({ S1965, S1801 }),
  .out1({ S1966 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2539_ (
  .in1({ S1966, S1857 }),
  .out1({ S1967 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2540_ (
  .in1({ S1856, S1754 }),
  .out1({ S1968 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2541_ (
  .in1({ S1968, S1967 }),
  .out1({ S1969 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2542_ (
  .in1({ S1969 }),
  .out1({ S1970 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2543_ (
  .in1({ S1970, S241 }),
  .out1({ S1971 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2544_ (
  .in1({ S1969, S240 }),
  .out1({ S1972 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2545_ (
  .in1({ S1969, S240 }),
  .out1({ S1973 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2546_ (
  .in1({ S1970, S241 }),
  .out1({ S1974 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2547_ (
  .in1({ S1796, S1775 }),
  .out1({ S1975 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2548_ (
  .in1({ S1975, S1797 }),
  .out1({ S1976 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2549_ (
  .in1({ S1976, S1857 }),
  .out1({ S1977 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2550_ (
  .in1({ S1977 }),
  .out1({ S1978 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2551_ (
  .in1({ S1856, S1769 }),
  .out1({ S1979 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2552_ (
  .in1({ S1857, S1770 }),
  .out1({ S1980 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2553_ (
  .in1({ S1979, S1977 }),
  .out1({ S1981 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2554_ (
  .in1({ S1980, S1978 }),
  .out1({ S1982 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2555_ (
  .in1({ S1982, S249 }),
  .out1({ S1983 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2556_ (
  .in1({ S1981, S248 }),
  .out1({ S1984 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2557_ (
  .in1({ S1981, S248 }),
  .out1({ S1985 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2558_ (
  .in1({ S1982, S249 }),
  .out1({ S1986 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2559_ (
  .in1({ S1985, S1983 }),
  .out1({ S1987 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2560_ (
  .in1({ S1986, S1984 }),
  .out1({ S1988 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2561_ (
  .in1({ S1791, S1788 }),
  .out1({ S1989 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2562_ (
  .in1({ S1989, S1793 }),
  .out1({ S1990 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2563_ (
  .in1({ S1990, S1857 }),
  .out1({ S1991 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2564_ (
  .in1({ S1991 }),
  .out1({ S1992 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2565_ (
  .in1({ S1856, S1784 }),
  .out1({ S1993 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2566_ (
  .in1({ S1857, S1783 }),
  .out1({ S1994 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2567_ (
  .in1({ S1993, S1991 }),
  .out1({ S1995 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2568_ (
  .in1({ S1994, S1992 }),
  .out1({ S1996 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2569_ (
  .in1({ S1996, S257 }),
  .out1({ S1997 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2570_ (
  .in1({ S1995, S256 }),
  .out1({ S1998 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2571_ (
  .in1({ S1995, S256 }),
  .out1({ S1999 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2572_ (
  .in1({ S1996, S257 }),
  .out1({ S2000 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2573_ (
  .in1({ S1999, S1997 }),
  .out1({ S2001 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2574_ (
  .in1({ S2000, S1998 }),
  .out1({ S2002 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2575_ (
  .in1({ S1857, S270 }),
  .out1({ S2003 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2576_ (
  .in1({ S1856, S271 }),
  .out1({ S2004 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2577_ (
  .in1({ S2004, S5957 }),
  .out1({ S2005 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2578_ (
  .in1({ S2003, new_datapath_addsubunit_in1_2 }),
  .out1({ S2006 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2579_ (
  .in1({ S2003, new_datapath_addsubunit_in1_2 }),
  .out1({ S2007 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2580_ (
  .in1({ S2004, S5957 }),
  .out1({ S2008 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2581_ (
  .in1({ S2008, S2006 }),
  .out1({ S2009 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2582_ (
  .in1({ S2007, S2005 }),
  .out1({ S2010 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2583_ (
  .in1({ S2009, S265 }),
  .out1({ S2011 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2584_ (
  .in1({ S2010, S264 }),
  .out1({ S2012 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2585_ (
  .in1({ S2010, S264 }),
  .out1({ S2013 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2586_ (
  .in1({ S2009, S265 }),
  .out1({ S2014 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2587_ (
  .in1({ S2013, S2011 }),
  .out1({ S2015 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2588_ (
  .in1({ S2014, S2012 }),
  .out1({ S2016 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2589_ (
  .in1({ S271, S5966 }),
  .out1({ S2017 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2590_ (
  .in1({ S2017 }),
  .out1({ S2018 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2591_ (
  .in1({ S2018, S2016 }),
  .out1({ S2019 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2592_ (
  .in1({ S2017, S2015 }),
  .out1({ S2020 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2593_ (
  .in1({ S2019, S2011 }),
  .out1({ S2021 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2594_ (
  .in1({ S2020, S2012 }),
  .out1({ S2022 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2595_ (
  .in1({ S2021, S2002 }),
  .out1({ S2023 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2596_ (
  .in1({ S2022, S2001 }),
  .out1({ S2024 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2597_ (
  .in1({ S2023, S1997 }),
  .out1({ S2025 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2598_ (
  .in1({ S2024, S1998 }),
  .out1({ S2026 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2599_ (
  .in1({ S2025, S1988 }),
  .out1({ S2027 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2600_ (
  .in1({ S2026, S1987 }),
  .out1({ S2028 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2601_ (
  .in1({ S2027, S1983 }),
  .out1({ S2029 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2602_ (
  .in1({ S2028, S1984 }),
  .out1({ S2030 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2603_ (
  .in1({ S2029, S1973 }),
  .out1({ S2031 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2604_ (
  .in1({ S2030, S1974 }),
  .out1({ S2032 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2605_ (
  .in1({ S2031, S1971 }),
  .out1({ S2033 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2606_ (
  .in1({ S2032, S1972 }),
  .out1({ S2034 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2607_ (
  .in1({ S2033, S1963 }),
  .out1({ S2035 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2608_ (
  .in1({ S2034, S1964 }),
  .out1({ S2036 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2609_ (
  .in1({ S2035, S1961 }),
  .out1({ S2037 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2610_ (
  .in1({ S2036, S1960 }),
  .out1({ S2038 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2611_ (
  .in1({ S2037, S1953 }),
  .out1({ S2039 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2612_ (
  .in1({ S2038, S1952 }),
  .out1({ S2040 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2613_ (
  .in1({ S2039, S1952 }),
  .out1({ S2041 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2614_ (
  .in1({ S2040, S1953 }),
  .out1({ S2042 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2615_ (
  .in1({ S2041, S1943 }),
  .out1({ S2043 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2616_ (
  .in1({ S2042, S1942 }),
  .out1({ S2044 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2617_ (
  .in1({ S2043, S1939 }),
  .out1({ S2045 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2618_ (
  .in1({ S2044, S1940 }),
  .out1({ S2046 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2619_ (
  .in1({ S2046, S1932 }),
  .out1({ S2047 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2620_ (
  .in1({ S2045, S1931 }),
  .out1({ S2048 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2621_ (
  .in1({ S2048, S1932 }),
  .out1({ S2049 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2622_ (
  .in1({ S2047, S1931 }),
  .out1({ S2050 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2623_ (
  .in1({ S2049, S1919 }),
  .out1({ S2051 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2624_ (
  .in1({ S2050, S1920 }),
  .out1({ S2052 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2625_ (
  .in1({ S2051, S1916 }),
  .out1({ S2053 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2626_ (
  .in1({ S2052, S1917 }),
  .out1({ S2054 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2627_ (
  .in1({ S2054, S1909 }),
  .out1({ S2055 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2628_ (
  .in1({ S2053, S1908 }),
  .out1({ S2056 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2629_ (
  .in1({ S2056, S1909 }),
  .out1({ S2057 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2630_ (
  .in1({ S2055, S1908 }),
  .out1({ S2058 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2631_ (
  .in1({ S2057, S1896 }),
  .out1({ S2059 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2632_ (
  .in1({ S2058, S1895 }),
  .out1({ S2060 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2633_ (
  .in1({ S2059, S1891 }),
  .out1({ S2061 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2634_ (
  .in1({ S2060, S1892 }),
  .out1({ S2062 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2635_ (
  .in1({ S2062, S1881 }),
  .out1({ S2063 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2636_ (
  .in1({ S2061, S1880 }),
  .out1({ S2064 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2637_ (
  .in1({ S2064, S1881 }),
  .out1({ S2065 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2638_ (
  .in1({ S2063, S1880 }),
  .out1({ S2066 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2639_ (
  .in1({ S2065, S1867 }),
  .out1({ S2067 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2640_ (
  .in1({ S2066, S1868 }),
  .out1({ S2068 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2641_ (
  .in1({ S2067, S1864 }),
  .out1({ S2069 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2642_ (
  .in1({ S2068, S1865 }),
  .out1({ S2070 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2643_ (
  .in1({ S210, new_datapath_multdivunit_1697_B_13 }),
  .out1({ S2071 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2644_ (
  .in1({ S2071, S1842 }),
  .out1({ S2072 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2645_ (
  .in1({ S1842, S212 }),
  .out1({ S2073 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2646_ (
  .in1({ S2072, S1848 }),
  .out1({ S2074 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2647_ (
  .in1({ S2074, S2073 }),
  .out1({ S2075 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2648_ (
  .in1({ S2075, new_datapath_multdivunit_1697_B_14 }),
  .out1({ S2076 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2649_ (
  .in1({ S2076 }),
  .out1({ S2077 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2650_ (
  .in1({ S2076, S2070 }),
  .out1({ S2078 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2651_ (
  .in1({ S2077, S2069 }),
  .out1({ S2079 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2652_ (
  .in1({ S2075, new_datapath_multdivunit_1697_B_15 }),
  .out1({ S2080 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2653_ (
  .in1({ S2080, S210 }),
  .out1({ S2081 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2654_ (
  .in1({ S2081 }),
  .out1({ S2082 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2655_ (
  .in1({ S2081, S2078 }),
  .out1({ S2083 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2656_ (
  .in1({ S2082, S2079 }),
  .out1({ S2084 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2657_ (
  .in1({ S2033, S1963 }),
  .out1({ S2085 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2658_ (
  .in1({ S2085, S2036 }),
  .out1({ S2086 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2659_ (
  .in1({ S2086, S2083 }),
  .out1({ S2087 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2660_ (
  .in1({ S2084, S1958 }),
  .out1({ S2088 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2661_ (
  .in1({ S2088, S2087 }),
  .out1({ S2089 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2662_ (
  .in1({ S2089, S203 }),
  .out1({ S2090 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2663_ (
  .in1({ S1973, S1971 }),
  .out1({ S2091 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2664_ (
  .in1({ S1974, S1972 }),
  .out1({ S2092 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2665_ (
  .in1({ S2091, S2029 }),
  .out1({ S2093 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2666_ (
  .in1({ S2092, S2030 }),
  .out1({ S2094 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2667_ (
  .in1({ S2094, S2093 }),
  .out1({ S2095 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2668_ (
  .in1({ S2095, S2084 }),
  .out1({ S2096 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2669_ (
  .in1({ S2083, S1969 }),
  .out1({ S2097 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2670_ (
  .in1({ S2097, S2096 }),
  .out1({ S2098 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2671_ (
  .in1({ S2098, S208 }),
  .out1({ S2099 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2672_ (
  .in1({ S2017, S2015 }),
  .out1({ S2100 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2673_ (
  .in1({ S2100, S2019 }),
  .out1({ S2101 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2674_ (
  .in1({ S2101, S2084 }),
  .out1({ S2102 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2675_ (
  .in1({ S2083, S2010 }),
  .out1({ S2103 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2676_ (
  .in1({ S2103, S2102 }),
  .out1({ S2104 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2677_ (
  .in1({ S2104, S256 }),
  .out1({ S2105 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2678_ (
  .in1({ S2083, S271 }),
  .out1({ S2106 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2679_ (
  .in1({ S2106, new_datapath_addsubunit_in1_1 }),
  .out1({ S2107 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2680_ (
  .in1({ S270, new_datapath_addsubunit_in1_0 }),
  .out1({ S2108 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2681_ (
  .in1({ S2108, S265 }),
  .out1({ S2109 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2682_ (
  .in1({ S2084, S2017 }),
  .out1({ S2110 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2683_ (
  .in1({ S2110, S2109 }),
  .out1({ S2111 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2684_ (
  .in1({ S2111, S2107 }),
  .out1({ S2112 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2685_ (
  .in1({ S2108, S265 }),
  .out1({ S2113 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2686_ (
  .in1({ S2113, S2112 }),
  .out1({ S2114 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2687_ (
  .in1({ S2114, S2105 }),
  .out1({ S2115 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2688_ (
  .in1({ S2083, S1995 }),
  .out1({ S2116 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2689_ (
  .in1({ S2084, S1996 }),
  .out1({ S2117 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2690_ (
  .in1({ S2022, S2001 }),
  .out1({ S2118 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2691_ (
  .in1({ S2021, S2002 }),
  .out1({ S2119 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2692_ (
  .in1({ S2118, S2023 }),
  .out1({ S2120 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2693_ (
  .in1({ S2119, S2024 }),
  .out1({ S2121 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2694_ (
  .in1({ S2120, S2084 }),
  .out1({ S2122 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2695_ (
  .in1({ S2121, S2083 }),
  .out1({ S2123 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2696_ (
  .in1({ S2122, S2116 }),
  .out1({ S2124 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2697_ (
  .in1({ S2123, S2117 }),
  .out1({ S2125 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2698_ (
  .in1({ S2124, S248 }),
  .out1({ S2126 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2699_ (
  .in1({ S2104, S256 }),
  .out1({ S2127 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2700_ (
  .in1({ S2127, S2126 }),
  .out1({ S2128 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2701_ (
  .in1({ S2128, S2115 }),
  .out1({ S2129 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2702_ (
  .in1({ S2125, S249 }),
  .out1({ S2130 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2703_ (
  .in1({ S2083, S1981 }),
  .out1({ S2131 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2704_ (
  .in1({ S2084, S1982 }),
  .out1({ S2132 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2705_ (
  .in1({ S2026, S1987 }),
  .out1({ S2133 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2706_ (
  .in1({ S2025, S1988 }),
  .out1({ S2134 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2707_ (
  .in1({ S2133, S2027 }),
  .out1({ S2135 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2708_ (
  .in1({ S2134, S2028 }),
  .out1({ S2136 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2709_ (
  .in1({ S2135, S2084 }),
  .out1({ S2137 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2710_ (
  .in1({ S2136, S2083 }),
  .out1({ S2138 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2711_ (
  .in1({ S2137, S2131 }),
  .out1({ S2139 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2712_ (
  .in1({ S2138, S2132 }),
  .out1({ S2140 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2713_ (
  .in1({ S2140, S241 }),
  .out1({ S2141 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2714_ (
  .in1({ S2141, S2130 }),
  .out1({ S2142 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2715_ (
  .in1({ S2142, S2129 }),
  .out1({ S2143 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2716_ (
  .in1({ S2098, S208 }),
  .out1({ S2144 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2717_ (
  .in1({ S2139, S240 }),
  .out1({ S2145 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2718_ (
  .in1({ S2145, S2144 }),
  .out1({ S2146 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2719_ (
  .in1({ S2146, S2143 }),
  .out1({ S2147 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2720_ (
  .in1({ S2147, S2099 }),
  .out1({ S2148 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2721_ (
  .in1({ S2148, S2090 }),
  .out1({ S2149 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2722_ (
  .in1({ S1953, S1952 }),
  .out1({ S2150 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2723_ (
  .in1({ S2150, S2038 }),
  .out1({ S2151 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2724_ (
  .in1({ S2151 }),
  .out1({ S2152 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2725_ (
  .in1({ S2150, S2038 }),
  .out1({ S2153 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2726_ (
  .in1({ S2153 }),
  .out1({ S2154 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2727_ (
  .in1({ S2154, S2151 }),
  .out1({ S2155 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2728_ (
  .in1({ S2153, S2152 }),
  .out1({ S2156 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2729_ (
  .in1({ S2155, S2084 }),
  .out1({ S2157 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2730_ (
  .in1({ S2156, S2083 }),
  .out1({ S2158 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2731_ (
  .in1({ S2083, S1950 }),
  .out1({ S2159 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2732_ (
  .in1({ S2084, S1951 }),
  .out1({ S2160 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2733_ (
  .in1({ S2159, S2157 }),
  .out1({ S2161 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2734_ (
  .in1({ S2160, S2158 }),
  .out1({ S2162 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2735_ (
  .in1({ S2162, S229 }),
  .out1({ S2163 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2736_ (
  .in1({ S2089, S203 }),
  .out1({ S2164 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2737_ (
  .in1({ S2164, S2163 }),
  .out1({ S2165 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2738_ (
  .in1({ S2165, S2149 }),
  .out1({ S2166 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2739_ (
  .in1({ S2083, S1907 }),
  .out1({ S2167 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2740_ (
  .in1({ S2084, S1906 }),
  .out1({ S2168 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2741_ (
  .in1({ S1909, S1908 }),
  .out1({ S2169 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2742_ (
  .in1({ S2169, S2053 }),
  .out1({ S2170 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2743_ (
  .in1({ S2170 }),
  .out1({ S2171 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2744_ (
  .in1({ S2169, S2053 }),
  .out1({ S2172 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2745_ (
  .in1({ S2172 }),
  .out1({ S2173 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2746_ (
  .in1({ S2172, S2171 }),
  .out1({ S2174 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2747_ (
  .in1({ S2173, S2170 }),
  .out1({ S2175 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2748_ (
  .in1({ S2175, S2084 }),
  .out1({ S2176 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2749_ (
  .in1({ S2174, S2083 }),
  .out1({ S2177 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2750_ (
  .in1({ S2176, S2167 }),
  .out1({ S2178 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2751_ (
  .in1({ S2177, S2168 }),
  .out1({ S2179 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2752_ (
  .in1({ S2178, new_datapath_multdivunit_1697_B_11 }),
  .out1({ S2180 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2753_ (
  .in1({ S2179, S3445 }),
  .out1({ S2181 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2754_ (
  .in1({ S2181, S2180 }),
  .out1({ S2182 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2755_ (
  .in1({ S2049, S1919 }),
  .out1({ S2183 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2756_ (
  .in1({ S2183, S2052 }),
  .out1({ S2184 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2757_ (
  .in1({ S2184, S2083 }),
  .out1({ S2185 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2758_ (
  .in1({ S2084, S1914 }),
  .out1({ S2186 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2759_ (
  .in1({ S2186, S2185 }),
  .out1({ S2187 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2760_ (
  .in1({ S2187, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S2188 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2761_ (
  .in1({ S2187, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S2189 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2762_ (
  .in1({ S2189 }),
  .out1({ S2190 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2763_ (
  .in1({ S2190, S2188 }),
  .out1({ S2191 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2764_ (
  .in1({ S2191, S2182 }),
  .out1({ S2192 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2765_ (
  .in1({ S2161, S228 }),
  .out1({ S2193 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2766_ (
  .in1({ S2042, S1942 }),
  .out1({ S2194 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2767_ (
  .in1({ S2194, S2043 }),
  .out1({ S2195 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2768_ (
  .in1({ S2195, S2084 }),
  .out1({ S2196 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2769_ (
  .in1({ S2083, S1937 }),
  .out1({ S2197 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2770_ (
  .in1({ S2197, S2196 }),
  .out1({ S2198 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2771_ (
  .in1({ S2198, S3478 }),
  .out1({ S2199 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2772_ (
  .in1({ S2199, S2193 }),
  .out1({ S2200 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2773_ (
  .in1({ S1932, S1931 }),
  .out1({ S2201 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2774_ (
  .in1({ S2201, S2045 }),
  .out1({ S2202 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2775_ (
  .in1({ S2202 }),
  .out1({ S2203 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2776_ (
  .in1({ S2201, S2045 }),
  .out1({ S2204 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2777_ (
  .in1({ S2204, S2203 }),
  .out1({ S2205 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2778_ (
  .in1({ S2205, S2084 }),
  .out1({ S2206 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2779_ (
  .in1({ S2083, S1929 }),
  .out1({ S2207 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2780_ (
  .in1({ S2207, S2206 }),
  .out1({ S2208 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2781_ (
  .in1({ S2208 }),
  .out1({ S2209 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2782_ (
  .in1({ S2208, S3467 }),
  .out1({ S2210 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2783_ (
  .in1({ S2209, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S2211 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2784_ (
  .in1({ S2208, S3467 }),
  .out1({ S2212 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2785_ (
  .in1({ S2198, S3478 }),
  .out1({ S2213 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2786_ (
  .in1({ S2213, S2212 }),
  .out1({ S2214 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2787_ (
  .in1({ S2214, S2210 }),
  .out1({ S2215 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2788_ (
  .in1({ S2215, S2200 }),
  .out1({ S2216 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2789_ (
  .in1({ S2216, S2192 }),
  .out1({ S2217 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2790_ (
  .in1({ S2217, S2166 }),
  .out1({ S2218 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2791_ (
  .in1({ S2214, S2211 }),
  .out1({ S2219 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2792_ (
  .in1({ S2219, S2192 }),
  .out1({ S2220 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2793_ (
  .in1({ S2188, S2180 }),
  .out1({ S2221 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2794_ (
  .in1({ S2221, S2181 }),
  .out1({ S2222 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2795_ (
  .in1({ S2222, S2220 }),
  .out1({ S2223 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2796_ (
  .in1({ S2223, S2218 }),
  .out1({ S2224 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2797_ (
  .in1({ S2065, S1867 }),
  .out1({ S2225 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2798_ (
  .in1({ S2225, S2068 }),
  .out1({ S2226 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2799_ (
  .in1({ S2226, S2083 }),
  .out1({ S2227 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2800_ (
  .in1({ S2084, S1862 }),
  .out1({ S2228 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2801_ (
  .in1({ S2228, S2227 }),
  .out1({ S2229 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2802_ (
  .in1({ S2069, S3412 }),
  .out1({ S2230 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2803_ (
  .in1({ S2230 }),
  .out1({ S2231 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2804_ (
  .in1({ S1848, new_datapath_multdivunit_1697_B_15 }),
  .out1({ S2232 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2805_ (
  .in1({ S2229, new_datapath_multdivunit_1697_B_14 }),
  .out1({ S2233 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2806_ (
  .in1({ S2233 }),
  .out1({ S2234 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2807_ (
  .in1({ S2229, new_datapath_multdivunit_1697_B_14 }),
  .out1({ S2235 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2808_ (
  .in1({ S2069, S3412 }),
  .out1({ S2236 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2809_ (
  .in1({ S2236, S2231 }),
  .out1({ S2237 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2810_ (
  .in1({ S2237, S2080 }),
  .out1({ S2238 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2811_ (
  .in1({ S2235, S2234 }),
  .out1({ S2239 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2812_ (
  .in1({ S2238, S2232 }),
  .out1({ S2240 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2813_ (
  .in1({ S2240 }),
  .out1({ S2241 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2814_ (
  .in1({ S2241, S2239 }),
  .out1({ S2242 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2815_ (
  .in1({ S1881, S1880 }),
  .out1({ S2243 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2816_ (
  .in1({ S2243, S2061 }),
  .out1({ S2244 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2817_ (
  .in1({ S2244 }),
  .out1({ S2245 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2818_ (
  .in1({ S2243, S2061 }),
  .out1({ S2246 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2819_ (
  .in1({ S2246 }),
  .out1({ S2247 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2820_ (
  .in1({ S2246, S2245 }),
  .out1({ S2248 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2821_ (
  .in1({ S2247, S2244 }),
  .out1({ S2249 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2822_ (
  .in1({ S2248, S2084 }),
  .out1({ S2250 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2823_ (
  .in1({ S2249, S2083 }),
  .out1({ S2251 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2824_ (
  .in1({ S2083, S1878 }),
  .out1({ S2252 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2825_ (
  .in1({ S2084, S1879 }),
  .out1({ S2253 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2826_ (
  .in1({ S2252, S2250 }),
  .out1({ S2254 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2827_ (
  .in1({ S2253, S2251 }),
  .out1({ S2255 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2828_ (
  .in1({ S2255, new_datapath_multdivunit_1697_B_13 }),
  .out1({ S2256 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2829_ (
  .in1({ S2254, S3423 }),
  .out1({ S2257 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2830_ (
  .in1({ S2058, S1895 }),
  .out1({ S2258 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2831_ (
  .in1({ S2258, S2059 }),
  .out1({ S2259 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2832_ (
  .in1({ S2259, S2084 }),
  .out1({ S2260 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2833_ (
  .in1({ S2083, S1889 }),
  .out1({ S2261 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2834_ (
  .in1({ S2261, S2260 }),
  .out1({ S2262 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2835_ (
  .in1({ S2262 }),
  .out1({ S2263 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2836_ (
  .in1({ S2263, new_datapath_multdivunit_1697_B_12 }),
  .out1({ S2264 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2837_ (
  .in1({ S2262, S3434 }),
  .out1({ S2265 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2838_ (
  .in1({ S2264, S2256 }),
  .out1({ S2266 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2839_ (
  .in1({ S2265, S2257 }),
  .out1({ S2267 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2840_ (
  .in1({ S2254, S3423 }),
  .out1({ S2268 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2841_ (
  .in1({ S2255, new_datapath_multdivunit_1697_B_13 }),
  .out1({ S2269 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2842_ (
  .in1({ S2262, S3434 }),
  .out1({ S2270 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2843_ (
  .in1({ S2270, S2268 }),
  .out1({ S2271 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2844_ (
  .in1({ S2271, S2266 }),
  .out1({ S2272 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2845_ (
  .in1({ S2272, S2242 }),
  .out1({ S2273 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2846_ (
  .in1({ S2273, S2224 }),
  .out1({ S2274 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2847_ (
  .in1({ S2269, S2267 }),
  .out1({ S2275 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2848_ (
  .in1({ S2275, S2242 }),
  .out1({ S2276 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2849_ (
  .in1({ S2235, S2232 }),
  .out1({ S2277 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2850_ (
  .in1({ S2277, S2238 }),
  .out1({ S2278 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2851_ (
  .in1({ S2278, S2276 }),
  .out1({ S2279 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2852_ (
  .in1({ S2279, S2274 }),
  .out1({ S2280 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2853_ (
  .in1({ S2280, S5537 }),
  .out1({ S2281 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2854_ (
  .in1({ S5611, new_datapath_multdivunit_outmdu1_0 }),
  .out1({ S2282 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2855_ (
  .in1({ S270, S5590 }),
  .out1({ S2283 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2856_ (
  .in1({ S2283, new_datapath_addsubunit_in1_0 }),
  .out1({ S2284 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2857_ (
  .in1({ S2284, S2282 }),
  .out1({ S2285 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2858_ (
  .in1({ S2285 }),
  .out1({ S2286 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2859_ (
  .in1({ S2286, S2281 }),
  .out1({ S20 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2860_ (
  .in1({ S2084, S5547 }),
  .out1({ S2287 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2861_ (
  .in1({ S5611, new_datapath_multdivunit_outmdu1_1 }),
  .out1({ S2288 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2862_ (
  .in1({ S270, S5966 }),
  .out1({ S2289 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2863_ (
  .in1({ S264, S5975 }),
  .out1({ S2290 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2864_ (
  .in1({ S265, new_datapath_addsubunit_in1_1 }),
  .out1({ S2291 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2865_ (
  .in1({ S2290, S2289 }),
  .out1({ S2292 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2866_ (
  .in1({ S2290, S2289 }),
  .out1({ S2293 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2867_ (
  .in1({ S2292, S5579 }),
  .out1({ S2294 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2868_ (
  .in1({ S2294, S2293 }),
  .out1({ S2295 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2869_ (
  .in1({ S2295, S2287 }),
  .out1({ S2296 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2870_ (
  .in1({ S2296, S2288 }),
  .out1({ S21 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2871_ (
  .in1({ S1857, S5547 }),
  .out1({ S2297 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2872_ (
  .in1({ S256, S5975 }),
  .out1({ S2298 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2873_ (
  .in1({ S257, new_datapath_addsubunit_in1_0 }),
  .out1({ S2299 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2874_ (
  .in1({ S271, new_datapath_addsubunit_in1_2 }),
  .out1({ S2300 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2875_ (
  .in1({ S2300, S2291 }),
  .out1({ S2301 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2876_ (
  .in1({ S264, S5957 }),
  .out1({ S2302 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2877_ (
  .in1({ S265, new_datapath_addsubunit_in1_2 }),
  .out1({ S2303 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2878_ (
  .in1({ S2302, S2289 }),
  .out1({ S2304 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2879_ (
  .in1({ S2304, S2301 }),
  .out1({ S2305 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2880_ (
  .in1({ S2305 }),
  .out1({ S2306 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2881_ (
  .in1({ S2306, S2298 }),
  .out1({ S2307 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2882_ (
  .in1({ S2305, S2299 }),
  .out1({ S2308 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2883_ (
  .in1({ S2308, S2307 }),
  .out1({ S2309 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2884_ (
  .in1({ S2309, S2292 }),
  .out1({ S2310 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2885_ (
  .in1({ S2309, S2292 }),
  .out1({ S2311 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2886_ (
  .in1({ S2311, S5590 }),
  .out1({ S2312 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2887_ (
  .in1({ S2312, S2310 }),
  .out1({ S2313 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2888_ (
  .in1({ S5611, new_datapath_multdivunit_outmdu1_2 }),
  .out1({ S2314 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2889_ (
  .in1({ S2314 }),
  .out1({ S2315 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2890_ (
  .in1({ S2315, S2297 }),
  .out1({ S2316 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2891_ (
  .in1({ S2316, S2313 }),
  .out1({ S22 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2892_ (
  .in1({ S1635, S5547 }),
  .out1({ S2317 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2893_ (
  .in1({ S5611, new_datapath_multdivunit_outmdu1_3 }),
  .out1({ S2318 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2894_ (
  .in1({ S248, S5975 }),
  .out1({ S2319 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2895_ (
  .in1({ S249, new_datapath_addsubunit_in1_0 }),
  .out1({ S2320 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2896_ (
  .in1({ S2307, S2304 }),
  .out1({ S2321 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2897_ (
  .in1({ S2321 }),
  .out1({ S2322 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2898_ (
  .in1({ S256, S5966 }),
  .out1({ S2323 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2899_ (
  .in1({ S257, new_datapath_addsubunit_in1_1 }),
  .out1({ S2324 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2900_ (
  .in1({ S270, S5947 }),
  .out1({ S2325 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2901_ (
  .in1({ S271, new_datapath_addsubunit_in1_3 }),
  .out1({ S2326 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2902_ (
  .in1({ S2325, S2302 }),
  .out1({ S2327 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2903_ (
  .in1({ S2326, S2303 }),
  .out1({ S2328 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2904_ (
  .in1({ S264, S5947 }),
  .out1({ S2329 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2905_ (
  .in1({ S265, new_datapath_addsubunit_in1_3 }),
  .out1({ S2330 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2906_ (
  .in1({ S2326, S2303 }),
  .out1({ S2331 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2907_ (
  .in1({ S2325, S2302 }),
  .out1({ S2332 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2908_ (
  .in1({ S2331, S2327 }),
  .out1({ S2333 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2909_ (
  .in1({ S2332, S2328 }),
  .out1({ S2334 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2910_ (
  .in1({ S2334, S2324 }),
  .out1({ S2335 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2911_ (
  .in1({ S2333, S2323 }),
  .out1({ S2336 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2912_ (
  .in1({ S2333, S2323 }),
  .out1({ S2337 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2913_ (
  .in1({ S2334, S2324 }),
  .out1({ S2338 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2914_ (
  .in1({ S2337, S2335 }),
  .out1({ S2339 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2915_ (
  .in1({ S2338, S2336 }),
  .out1({ S2340 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2916_ (
  .in1({ S2340, S2322 }),
  .out1({ S2341 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2917_ (
  .in1({ S2339, S2321 }),
  .out1({ S2342 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2918_ (
  .in1({ S2342, S2341 }),
  .out1({ S2343 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2919_ (
  .in1({ S2343 }),
  .out1({ S2344 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2920_ (
  .in1({ S2344, S2320 }),
  .out1({ S2345 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2921_ (
  .in1({ S2343, S2319 }),
  .out1({ S2346 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2922_ (
  .in1({ S2346, S2345 }),
  .out1({ S2347 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2923_ (
  .in1({ S2347, S2311 }),
  .out1({ S2348 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2924_ (
  .in1({ S2347, S2311 }),
  .out1({ S2349 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2925_ (
  .in1({ S2348, S5579 }),
  .out1({ S2350 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2926_ (
  .in1({ S2350, S2349 }),
  .out1({ S2351 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2927_ (
  .in1({ S2351, S2317 }),
  .out1({ S2352 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2928_ (
  .in1({ S2352, S2318 }),
  .out1({ S23 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2929_ (
  .in1({ S1452, S5547 }),
  .out1({ S2353 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2930_ (
  .in1({ S5611, new_datapath_multdivunit_outmdu1_4 }),
  .out1({ S2354 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2931_ (
  .in1({ S2345, S2341 }),
  .out1({ S2355 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2932_ (
  .in1({ S2355 }),
  .out1({ S2356 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2933_ (
  .in1({ S241, new_datapath_addsubunit_in1_0 }),
  .out1({ S2357 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2934_ (
  .in1({ S249, new_datapath_addsubunit_in1_1 }),
  .out1({ S2358 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2935_ (
  .in1({ S2358, S2357 }),
  .out1({ S2359 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2936_ (
  .in1({ S240, S5966 }),
  .out1({ S2360 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2937_ (
  .in1({ S241, new_datapath_addsubunit_in1_1 }),
  .out1({ S2361 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2938_ (
  .in1({ S2361, S2320 }),
  .out1({ S2362 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2939_ (
  .in1({ S2360, S2319 }),
  .out1({ S2363 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2940_ (
  .in1({ S2363, S2359 }),
  .out1({ S2364 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2941_ (
  .in1({ S2364 }),
  .out1({ S2365 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2942_ (
  .in1({ S2335, S2331 }),
  .out1({ S2366 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2943_ (
  .in1({ S2336, S2332 }),
  .out1({ S2367 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2944_ (
  .in1({ S256, S5957 }),
  .out1({ S2368 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2945_ (
  .in1({ S257, new_datapath_addsubunit_in1_2 }),
  .out1({ S2369 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2946_ (
  .in1({ S2329, S1204 }),
  .out1({ S2370 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2947_ (
  .in1({ S2330, S1205 }),
  .out1({ S2371 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2948_ (
  .in1({ S264, S5936 }),
  .out1({ S2372 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2949_ (
  .in1({ S265, new_datapath_addsubunit_in1_4 }),
  .out1({ S2373 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2950_ (
  .in1({ S2330, S1205 }),
  .out1({ S2374 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2951_ (
  .in1({ S2329, S1204 }),
  .out1({ S2375 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2952_ (
  .in1({ S2374, S2370 }),
  .out1({ S2376 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2953_ (
  .in1({ S2375, S2371 }),
  .out1({ S2377 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2954_ (
  .in1({ S2377, S2369 }),
  .out1({ S2378 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2955_ (
  .in1({ S2376, S2368 }),
  .out1({ S2379 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2956_ (
  .in1({ S2376, S2368 }),
  .out1({ S2380 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2957_ (
  .in1({ S2377, S2369 }),
  .out1({ S2381 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2958_ (
  .in1({ S2380, S2378 }),
  .out1({ S2382 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2959_ (
  .in1({ S2381, S2379 }),
  .out1({ S2383 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2960_ (
  .in1({ S2383, S2366 }),
  .out1({ S2384 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2961_ (
  .in1({ S2382, S2367 }),
  .out1({ S2385 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2962_ (
  .in1({ S2383, S2366 }),
  .out1({ S2386 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2963_ (
  .in1({ S2386, S2385 }),
  .out1({ S2387 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2964_ (
  .in1({ S2387 }),
  .out1({ S2388 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2965_ (
  .in1({ S2388, S2365 }),
  .out1({ S2389 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2966_ (
  .in1({ S2389 }),
  .out1({ S2390 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2967_ (
  .in1({ S2387, S2364 }),
  .out1({ S2391 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2968_ (
  .in1({ S2391, S2389 }),
  .out1({ S2392 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2969_ (
  .in1({ S2392 }),
  .out1({ S2393 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2970_ (
  .in1({ S2392, S2355 }),
  .out1({ S2394 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2971_ (
  .in1({ S2393, S2356 }),
  .out1({ S2395 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2972_ (
  .in1({ S2395 }),
  .out1({ S2396 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2973_ (
  .in1({ S2395, S2394 }),
  .out1({ S2397 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2974_ (
  .in1({ S2397, S2348 }),
  .out1({ S2398 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_2975_ (
  .in1({ S2398 }),
  .out1({ S2399 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2976_ (
  .in1({ S2397, S2348 }),
  .out1({ S2400 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2977_ (
  .in1({ S2400, S5579 }),
  .out1({ S2401 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2978_ (
  .in1({ S2401, S2398 }),
  .out1({ S2402 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2979_ (
  .in1({ S2402, S2353 }),
  .out1({ S2403 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2980_ (
  .in1({ S2403, S2354 }),
  .out1({ S24 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2981_ (
  .in1({ S1267, S5537 }),
  .out1({ S2404 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2982_ (
  .in1({ S2390, S2384 }),
  .out1({ S2405 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2983_ (
  .in1({ S2389, S2385 }),
  .out1({ S2406 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2984_ (
  .in1({ S208, S5975 }),
  .out1({ S2407 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2985_ (
  .in1({ S209, new_datapath_addsubunit_in1_0 }),
  .out1({ S2408 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2986_ (
  .in1({ S248, S5957 }),
  .out1({ S2409 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2987_ (
  .in1({ S249, new_datapath_addsubunit_in1_2 }),
  .out1({ S2410 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2988_ (
  .in1({ S2409, S2360 }),
  .out1({ S2411 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2989_ (
  .in1({ S2410, S2361 }),
  .out1({ S2412 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2990_ (
  .in1({ S240, S5957 }),
  .out1({ S2413 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2991_ (
  .in1({ S241, new_datapath_addsubunit_in1_2 }),
  .out1({ S2414 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2992_ (
  .in1({ S2410, S2361 }),
  .out1({ S2415 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2993_ (
  .in1({ S2409, S2360 }),
  .out1({ S2416 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2994_ (
  .in1({ S2415, S2411 }),
  .out1({ S2417 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2995_ (
  .in1({ S2416, S2412 }),
  .out1({ S2418 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2996_ (
  .in1({ S2418, S2408 }),
  .out1({ S2419 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2997_ (
  .in1({ S2417, S2407 }),
  .out1({ S2420 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_2998_ (
  .in1({ S2417, S2407 }),
  .out1({ S2421 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_2999_ (
  .in1({ S2418, S2408 }),
  .out1({ S2422 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3000_ (
  .in1({ S2421, S2419 }),
  .out1({ S2423 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3001_ (
  .in1({ S2422, S2420 }),
  .out1({ S2424 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3002_ (
  .in1({ S2378, S2374 }),
  .out1({ S2425 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3003_ (
  .in1({ S2379, S2375 }),
  .out1({ S2426 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3004_ (
  .in1({ S256, S5947 }),
  .out1({ S2427 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3005_ (
  .in1({ S257, new_datapath_addsubunit_in1_3 }),
  .out1({ S2428 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3006_ (
  .in1({ S2372, S1208 }),
  .out1({ S2429 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3007_ (
  .in1({ S2373, S1209 }),
  .out1({ S2430 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3008_ (
  .in1({ S264, S5926 }),
  .out1({ S2431 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3009_ (
  .in1({ S265, new_datapath_addsubunit_in1_5 }),
  .out1({ S2432 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3010_ (
  .in1({ S2373, S1209 }),
  .out1({ S2433 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3011_ (
  .in1({ S2372, S1208 }),
  .out1({ S2434 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3012_ (
  .in1({ S2433, S2429 }),
  .out1({ S2435 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3013_ (
  .in1({ S2434, S2430 }),
  .out1({ S2436 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3014_ (
  .in1({ S2436, S2428 }),
  .out1({ S2437 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3015_ (
  .in1({ S2435, S2427 }),
  .out1({ S2438 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3016_ (
  .in1({ S2435, S2427 }),
  .out1({ S2439 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3017_ (
  .in1({ S2436, S2428 }),
  .out1({ S2440 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3018_ (
  .in1({ S2439, S2437 }),
  .out1({ S2441 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3019_ (
  .in1({ S2440, S2438 }),
  .out1({ S2442 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3020_ (
  .in1({ S2442, S2425 }),
  .out1({ S2443 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3021_ (
  .in1({ S2441, S2426 }),
  .out1({ S2444 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3022_ (
  .in1({ S2441, S2426 }),
  .out1({ S2445 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3023_ (
  .in1({ S2442, S2425 }),
  .out1({ S2446 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3024_ (
  .in1({ S2445, S2443 }),
  .out1({ S2447 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3025_ (
  .in1({ S2446, S2444 }),
  .out1({ S2448 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3026_ (
  .in1({ S2448, S2424 }),
  .out1({ S2449 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3027_ (
  .in1({ S2447, S2423 }),
  .out1({ S2450 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3028_ (
  .in1({ S2447, S2423 }),
  .out1({ S2451 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3029_ (
  .in1({ S2448, S2424 }),
  .out1({ S2452 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3030_ (
  .in1({ S2451, S2449 }),
  .out1({ S2453 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3031_ (
  .in1({ S2452, S2450 }),
  .out1({ S2454 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3032_ (
  .in1({ S2453, S2406 }),
  .out1({ S2455 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3033_ (
  .in1({ S2454, S2405 }),
  .out1({ S2456 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3034_ (
  .in1({ S2456, S2455 }),
  .out1({ S2457 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3035_ (
  .in1({ S2457 }),
  .out1({ S2458 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3036_ (
  .in1({ S2458, S2362 }),
  .out1({ S2459 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3037_ (
  .in1({ S2457, S2363 }),
  .out1({ S2460 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3038_ (
  .in1({ S2460, S2459 }),
  .out1({ S2461 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3039_ (
  .in1({ S2461 }),
  .out1({ S2462 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3040_ (
  .in1({ S2462, S2396 }),
  .out1({ S2463 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3041_ (
  .in1({ S2461, S2395 }),
  .out1({ S2464 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3042_ (
  .in1({ S2464, S2463 }),
  .out1({ S2465 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3043_ (
  .in1({ S2465, S2399 }),
  .out1({ S2466 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3044_ (
  .in1({ S2466 }),
  .out1({ S2467 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3045_ (
  .in1({ S2465, S2399 }),
  .out1({ S2468 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3046_ (
  .in1({ S2468, S5579 }),
  .out1({ S2469 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3047_ (
  .in1({ S2469, S2466 }),
  .out1({ S2470 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3048_ (
  .in1({ S5611, new_datapath_multdivunit_outmdu1_5 }),
  .out1({ S2471 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3049_ (
  .in1({ S2471 }),
  .out1({ S2472 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3050_ (
  .in1({ S2472, S2470 }),
  .out1({ S2473 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3051_ (
  .in1({ S2473, S2404 }),
  .out1({ S25 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3052_ (
  .in1({ S1084, S5537 }),
  .out1({ S2474 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3053_ (
  .in1({ S5600, S2789 }),
  .out1({ S2475 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3054_ (
  .in1({ S2459, S2455 }),
  .out1({ S2476 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3055_ (
  .in1({ S2476 }),
  .out1({ S2477 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3056_ (
  .in1({ S202, S5975 }),
  .out1({ S2478 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3057_ (
  .in1({ S203, new_datapath_addsubunit_in1_0 }),
  .out1({ S2479 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3058_ (
  .in1({ S2419, S2415 }),
  .out1({ S2480 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3059_ (
  .in1({ S2420, S2416 }),
  .out1({ S2481 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3060_ (
  .in1({ S2480, S2479 }),
  .out1({ S2482 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3061_ (
  .in1({ S2481, S2478 }),
  .out1({ S2483 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3062_ (
  .in1({ S2481, S2478 }),
  .out1({ S2484 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3063_ (
  .in1({ S2480, S2479 }),
  .out1({ S2485 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3064_ (
  .in1({ S2484, S2482 }),
  .out1({ S2486 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3065_ (
  .in1({ S2485, S2483 }),
  .out1({ S2487 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3066_ (
  .in1({ S2449, S2443 }),
  .out1({ S2488 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3067_ (
  .in1({ S2450, S2444 }),
  .out1({ S2489 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3068_ (
  .in1({ S208, S5966 }),
  .out1({ S2490 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3069_ (
  .in1({ S209, new_datapath_addsubunit_in1_1 }),
  .out1({ S2491 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3070_ (
  .in1({ S248, S5947 }),
  .out1({ S2492 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3071_ (
  .in1({ S249, new_datapath_addsubunit_in1_3 }),
  .out1({ S2493 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3072_ (
  .in1({ S2492, S2413 }),
  .out1({ S2494 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3073_ (
  .in1({ S2493, S2414 }),
  .out1({ S2495 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3074_ (
  .in1({ S240, S5947 }),
  .out1({ S2496 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3075_ (
  .in1({ S241, new_datapath_addsubunit_in1_3 }),
  .out1({ S2497 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3076_ (
  .in1({ S2493, S2414 }),
  .out1({ S2498 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3077_ (
  .in1({ S2492, S2413 }),
  .out1({ S2499 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3078_ (
  .in1({ S2498, S2494 }),
  .out1({ S2500 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3079_ (
  .in1({ S2499, S2495 }),
  .out1({ S2501 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3080_ (
  .in1({ S2501, S2491 }),
  .out1({ S2502 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3081_ (
  .in1({ S2500, S2490 }),
  .out1({ S2503 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3082_ (
  .in1({ S2500, S2490 }),
  .out1({ S2504 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3083_ (
  .in1({ S2501, S2491 }),
  .out1({ S2505 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3084_ (
  .in1({ S2504, S2502 }),
  .out1({ S2506 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3085_ (
  .in1({ S2505, S2503 }),
  .out1({ S2507 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3086_ (
  .in1({ S2437, S2433 }),
  .out1({ S2508 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3087_ (
  .in1({ S2438, S2434 }),
  .out1({ S2509 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3088_ (
  .in1({ S256, S5936 }),
  .out1({ S2510 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3089_ (
  .in1({ S257, new_datapath_addsubunit_in1_4 }),
  .out1({ S2511 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3090_ (
  .in1({ S2431, S882 }),
  .out1({ S2512 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3091_ (
  .in1({ S2432, S883 }),
  .out1({ S2513 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3092_ (
  .in1({ S264, S5916 }),
  .out1({ S2514 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3093_ (
  .in1({ S265, new_datapath_addsubunit_in1_6 }),
  .out1({ S2515 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3094_ (
  .in1({ S2432, S883 }),
  .out1({ S2516 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3095_ (
  .in1({ S2431, S882 }),
  .out1({ S2517 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3096_ (
  .in1({ S2516, S2512 }),
  .out1({ S2518 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3097_ (
  .in1({ S2517, S2513 }),
  .out1({ S2519 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3098_ (
  .in1({ S2519, S2511 }),
  .out1({ S2520 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3099_ (
  .in1({ S2518, S2510 }),
  .out1({ S2521 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3100_ (
  .in1({ S2518, S2510 }),
  .out1({ S2522 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3101_ (
  .in1({ S2519, S2511 }),
  .out1({ S2523 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3102_ (
  .in1({ S2522, S2520 }),
  .out1({ S2524 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3103_ (
  .in1({ S2523, S2521 }),
  .out1({ S2525 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3104_ (
  .in1({ S2525, S2508 }),
  .out1({ S2526 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3105_ (
  .in1({ S2524, S2509 }),
  .out1({ S2527 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3106_ (
  .in1({ S2524, S2509 }),
  .out1({ S2528 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3107_ (
  .in1({ S2525, S2508 }),
  .out1({ S2529 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3108_ (
  .in1({ S2528, S2526 }),
  .out1({ S2530 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3109_ (
  .in1({ S2529, S2527 }),
  .out1({ S2531 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3110_ (
  .in1({ S2531, S2507 }),
  .out1({ S2532 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3111_ (
  .in1({ S2530, S2506 }),
  .out1({ S2533 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3112_ (
  .in1({ S2530, S2506 }),
  .out1({ S2534 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3113_ (
  .in1({ S2531, S2507 }),
  .out1({ S2535 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3114_ (
  .in1({ S2534, S2532 }),
  .out1({ S2536 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3115_ (
  .in1({ S2535, S2533 }),
  .out1({ S2537 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3116_ (
  .in1({ S2537, S2488 }),
  .out1({ S2538 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3117_ (
  .in1({ S2536, S2489 }),
  .out1({ S2539 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3118_ (
  .in1({ S2536, S2489 }),
  .out1({ S2540 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3119_ (
  .in1({ S2537, S2488 }),
  .out1({ S2541 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3120_ (
  .in1({ S2540, S2538 }),
  .out1({ S2542 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3121_ (
  .in1({ S2541, S2539 }),
  .out1({ S2543 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3122_ (
  .in1({ S2543, S2487 }),
  .out1({ S2544 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3123_ (
  .in1({ S2542, S2486 }),
  .out1({ S2545 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3124_ (
  .in1({ S2542, S2486 }),
  .out1({ S2546 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3125_ (
  .in1({ S2543, S2487 }),
  .out1({ S2547 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3126_ (
  .in1({ S2546, S2544 }),
  .out1({ S2548 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3127_ (
  .in1({ S2547, S2545 }),
  .out1({ S2549 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3128_ (
  .in1({ S2549, S2477 }),
  .out1({ S2550 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3129_ (
  .in1({ S2548, S2476 }),
  .out1({ S2551 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3130_ (
  .in1({ S2551 }),
  .out1({ S2552 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3131_ (
  .in1({ S2551, S2550 }),
  .out1({ S2553 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3132_ (
  .in1({ S2553, S2463 }),
  .out1({ S2554 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3133_ (
  .in1({ S2553, S2463 }),
  .out1({ S2555 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3134_ (
  .in1({ S2555 }),
  .out1({ S2556 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3135_ (
  .in1({ S2556, S2554 }),
  .out1({ S2557 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3136_ (
  .in1({ S2557 }),
  .out1({ S2558 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3137_ (
  .in1({ S2558, S2467 }),
  .out1({ S2559 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3138_ (
  .in1({ S2558, S2467 }),
  .out1({ S2560 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3139_ (
  .in1({ S2560, S5579 }),
  .out1({ S2561 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3140_ (
  .in1({ S2561, S2559 }),
  .out1({ S2562 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3141_ (
  .in1({ S2562, S2475 }),
  .out1({ S2563 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3142_ (
  .in1({ S2563, S2474 }),
  .out1({ S26 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3143_ (
  .in1({ S937, S5547 }),
  .out1({ S2564 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3144_ (
  .in1({ S5611, new_datapath_multdivunit_outmdu1_7 }),
  .out1({ S2565 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3145_ (
  .in1({ S2544, S2538 }),
  .out1({ S2566 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3146_ (
  .in1({ S2545, S2539 }),
  .out1({ S2567 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3147_ (
  .in1({ S228, S5975 }),
  .out1({ S2568 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3148_ (
  .in1({ S229, new_datapath_addsubunit_in1_0 }),
  .out1({ S2569 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3149_ (
  .in1({ S202, S5966 }),
  .out1({ S2570 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3150_ (
  .in1({ S203, new_datapath_addsubunit_in1_1 }),
  .out1({ S2571 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3151_ (
  .in1({ S2570, S2568 }),
  .out1({ S2572 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3152_ (
  .in1({ S2571, S2569 }),
  .out1({ S2573 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3153_ (
  .in1({ S228, S5966 }),
  .out1({ S2574 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3154_ (
  .in1({ S229, new_datapath_addsubunit_in1_1 }),
  .out1({ S2575 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3155_ (
  .in1({ S2575, S2479 }),
  .out1({ S2576 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3156_ (
  .in1({ S2574, S2478 }),
  .out1({ S2577 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3157_ (
  .in1({ S2576, S2572 }),
  .out1({ S2578 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3158_ (
  .in1({ S2577, S2573 }),
  .out1({ S2579 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3159_ (
  .in1({ S2502, S2498 }),
  .out1({ S2580 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3160_ (
  .in1({ S2503, S2499 }),
  .out1({ S2582 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3161_ (
  .in1({ S2582, S2578 }),
  .out1({ S2583 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3162_ (
  .in1({ S2580, S2579 }),
  .out1({ S2584 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3163_ (
  .in1({ S2580, S2579 }),
  .out1({ S2585 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3164_ (
  .in1({ S2582, S2578 }),
  .out1({ S2586 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3165_ (
  .in1({ S2585, S2583 }),
  .out1({ S2587 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3166_ (
  .in1({ S2586, S2584 }),
  .out1({ S2588 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3167_ (
  .in1({ S2532, S2526 }),
  .out1({ S2589 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3168_ (
  .in1({ S2533, S2527 }),
  .out1({ S2590 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3169_ (
  .in1({ S208, S5957 }),
  .out1({ S2591 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3170_ (
  .in1({ S209, new_datapath_addsubunit_in1_2 }),
  .out1({ S2593 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3171_ (
  .in1({ S248, S5936 }),
  .out1({ S2594 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3172_ (
  .in1({ S249, new_datapath_addsubunit_in1_4 }),
  .out1({ S2595 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3173_ (
  .in1({ S2594, S2496 }),
  .out1({ S2596 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3174_ (
  .in1({ S2595, S2497 }),
  .out1({ S2597 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3175_ (
  .in1({ S240, S5936 }),
  .out1({ S2598 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3176_ (
  .in1({ S241, new_datapath_addsubunit_in1_4 }),
  .out1({ S2599 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3177_ (
  .in1({ S2595, S2497 }),
  .out1({ S2600 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3178_ (
  .in1({ S2594, S2496 }),
  .out1({ S2601 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3179_ (
  .in1({ S2600, S2596 }),
  .out1({ S2602 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3180_ (
  .in1({ S2601, S2597 }),
  .out1({ S2604 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3181_ (
  .in1({ S2604, S2593 }),
  .out1({ S2605 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3182_ (
  .in1({ S2602, S2591 }),
  .out1({ S2606 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3183_ (
  .in1({ S2602, S2591 }),
  .out1({ S2607 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3184_ (
  .in1({ S2604, S2593 }),
  .out1({ S2608 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3185_ (
  .in1({ S2607, S2605 }),
  .out1({ S2609 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3186_ (
  .in1({ S2608, S2606 }),
  .out1({ S2610 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3187_ (
  .in1({ S2520, S2516 }),
  .out1({ S2611 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3188_ (
  .in1({ S2521, S2517 }),
  .out1({ S2612 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3189_ (
  .in1({ S256, S5926 }),
  .out1({ S2613 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3190_ (
  .in1({ S257, new_datapath_addsubunit_in1_5 }),
  .out1({ S2615 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3191_ (
  .in1({ S2514, S886 }),
  .out1({ S2616 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3192_ (
  .in1({ S2515, S887 }),
  .out1({ S2617 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3193_ (
  .in1({ S265, new_datapath_addsubunit_in1_7 }),
  .out1({ S2618 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3194_ (
  .in1({ S2515, S887 }),
  .out1({ S2619 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3195_ (
  .in1({ S2514, S886 }),
  .out1({ S2620 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3196_ (
  .in1({ S2619, S2616 }),
  .out1({ S2621 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3197_ (
  .in1({ S2620, S2617 }),
  .out1({ S2622 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3198_ (
  .in1({ S2622, S2615 }),
  .out1({ S2623 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3199_ (
  .in1({ S2621, S2613 }),
  .out1({ S2624 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3200_ (
  .in1({ S2621, S2613 }),
  .out1({ S2626 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3201_ (
  .in1({ S2622, S2615 }),
  .out1({ S2627 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3202_ (
  .in1({ S2626, S2623 }),
  .out1({ S2628 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3203_ (
  .in1({ S2627, S2624 }),
  .out1({ S2629 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3204_ (
  .in1({ S2629, S2611 }),
  .out1({ S2630 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3205_ (
  .in1({ S2628, S2612 }),
  .out1({ S2631 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3206_ (
  .in1({ S2628, S2612 }),
  .out1({ S2632 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3207_ (
  .in1({ S2629, S2611 }),
  .out1({ S2633 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3208_ (
  .in1({ S2632, S2630 }),
  .out1({ S2634 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3209_ (
  .in1({ S2633, S2631 }),
  .out1({ S2635 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3210_ (
  .in1({ S2635, S2610 }),
  .out1({ S2637 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3211_ (
  .in1({ S2634, S2609 }),
  .out1({ S2638 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3212_ (
  .in1({ S2634, S2609 }),
  .out1({ S2639 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3213_ (
  .in1({ S2635, S2610 }),
  .out1({ S2640 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3214_ (
  .in1({ S2639, S2637 }),
  .out1({ S2641 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3215_ (
  .in1({ S2640, S2638 }),
  .out1({ S2642 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3216_ (
  .in1({ S2642, S2589 }),
  .out1({ S2643 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3217_ (
  .in1({ S2641, S2590 }),
  .out1({ S2644 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3218_ (
  .in1({ S2641, S2590 }),
  .out1({ S2645 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3219_ (
  .in1({ S2642, S2589 }),
  .out1({ S2646 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3220_ (
  .in1({ S2645, S2643 }),
  .out1({ S2648 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3221_ (
  .in1({ S2646, S2644 }),
  .out1({ S2649 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3222_ (
  .in1({ S2649, S2588 }),
  .out1({ S2650 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3223_ (
  .in1({ S2648, S2587 }),
  .out1({ S2651 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3224_ (
  .in1({ S2648, S2587 }),
  .out1({ S2652 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3225_ (
  .in1({ S2649, S2588 }),
  .out1({ S2653 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3226_ (
  .in1({ S2652, S2650 }),
  .out1({ S2654 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3227_ (
  .in1({ S2653, S2651 }),
  .out1({ S2655 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3228_ (
  .in1({ S2655, S2566 }),
  .out1({ S2656 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3229_ (
  .in1({ S2654, S2567 }),
  .out1({ S2657 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3230_ (
  .in1({ S2655, S2566 }),
  .out1({ S2659 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3231_ (
  .in1({ S2659, S2657 }),
  .out1({ S2660 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3232_ (
  .in1({ S2660 }),
  .out1({ S2661 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3233_ (
  .in1({ S2661, S2482 }),
  .out1({ S2662 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3234_ (
  .in1({ S2662 }),
  .out1({ S2663 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3235_ (
  .in1({ S2660, S2483 }),
  .out1({ S2664 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3236_ (
  .in1({ S2664, S2662 }),
  .out1({ S2665 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3237_ (
  .in1({ S2665 }),
  .out1({ S2666 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3238_ (
  .in1({ S2666, S2552 }),
  .out1({ S2667 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3239_ (
  .in1({ S2667 }),
  .out1({ S2668 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3240_ (
  .in1({ S2665, S2551 }),
  .out1({ S2670 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3241_ (
  .in1({ S2670, S2667 }),
  .out1({ S2671 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3242_ (
  .in1({ S2671 }),
  .out1({ S2672 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3243_ (
  .in1({ S2672, S2559 }),
  .out1({ S2673 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3244_ (
  .in1({ S2673, S5579 }),
  .out1({ S2674 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3245_ (
  .in1({ S2559, S2554 }),
  .out1({ S2675 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3246_ (
  .in1({ S2675, S2671 }),
  .out1({ S2676 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3247_ (
  .in1({ S2672, S2554 }),
  .out1({ S2677 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3248_ (
  .in1({ S2677, S2676 }),
  .out1({ S2678 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3249_ (
  .in1({ S2678, S2674 }),
  .out1({ S2679 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3250_ (
  .in1({ S2679, S2564 }),
  .out1({ S2681 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3251_ (
  .in1({ S2681, S2565 }),
  .out1({ S27 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3252_ (
  .in1({ S788, S5547 }),
  .out1({ S2682 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3253_ (
  .in1({ S5611, new_datapath_multdivunit_outmdu1_8 }),
  .out1({ S2683 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3254_ (
  .in1({ S2663, S2656 }),
  .out1({ S2684 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3255_ (
  .in1({ S2662, S2657 }),
  .out1({ S2685 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3256_ (
  .in1({ S2650, S2643 }),
  .out1({ S2686 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3257_ (
  .in1({ S2651, S2644 }),
  .out1({ S2687 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3258_ (
  .in1({ S5975, S3478 }),
  .out1({ S2688 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3259_ (
  .in1({ new_datapath_addsubunit_in1_0, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S2689 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3260_ (
  .in1({ S202, S5957 }),
  .out1({ S2691 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3261_ (
  .in1({ S203, new_datapath_addsubunit_in1_2 }),
  .out1({ S2692 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3262_ (
  .in1({ S2691, S2574 }),
  .out1({ S2693 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3263_ (
  .in1({ S2692, S2575 }),
  .out1({ S2694 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3264_ (
  .in1({ S228, S5957 }),
  .out1({ S2695 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3265_ (
  .in1({ S229, new_datapath_addsubunit_in1_2 }),
  .out1({ S2696 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3266_ (
  .in1({ S2692, S2575 }),
  .out1({ S2697 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3267_ (
  .in1({ S2691, S2574 }),
  .out1({ S2698 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3268_ (
  .in1({ S2697, S2693 }),
  .out1({ S2699 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3269_ (
  .in1({ S2698, S2694 }),
  .out1({ S2700 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3270_ (
  .in1({ S2700, S2689 }),
  .out1({ S2702 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3271_ (
  .in1({ S2699, S2688 }),
  .out1({ S2703 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3272_ (
  .in1({ S2699, S2688 }),
  .out1({ S2704 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3273_ (
  .in1({ S2700, S2689 }),
  .out1({ S2705 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3274_ (
  .in1({ S2704, S2702 }),
  .out1({ S2706 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3275_ (
  .in1({ S2705, S2703 }),
  .out1({ S2707 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3276_ (
  .in1({ S2605, S2600 }),
  .out1({ S2708 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3277_ (
  .in1({ S2606, S2601 }),
  .out1({ S2709 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3278_ (
  .in1({ S2708, S2707 }),
  .out1({ S2710 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3279_ (
  .in1({ S2709, S2706 }),
  .out1({ S2711 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3280_ (
  .in1({ S2709, S2706 }),
  .out1({ S2713 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3281_ (
  .in1({ S2708, S2707 }),
  .out1({ S2714 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3282_ (
  .in1({ S2713, S2710 }),
  .out1({ S2715 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3283_ (
  .in1({ S2714, S2711 }),
  .out1({ S2716 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3284_ (
  .in1({ S2716, S2577 }),
  .out1({ S2717 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3285_ (
  .in1({ S2715, S2576 }),
  .out1({ S2718 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3286_ (
  .in1({ S2715, S2576 }),
  .out1({ S2719 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3287_ (
  .in1({ S2716, S2577 }),
  .out1({ S2720 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3288_ (
  .in1({ S2719, S2717 }),
  .out1({ S2721 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3289_ (
  .in1({ S2720, S2718 }),
  .out1({ S2722 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3290_ (
  .in1({ S2637, S2630 }),
  .out1({ S2724 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3291_ (
  .in1({ S2638, S2631 }),
  .out1({ S2725 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3292_ (
  .in1({ S208, S5947 }),
  .out1({ S2726 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3293_ (
  .in1({ S209, new_datapath_addsubunit_in1_3 }),
  .out1({ S2727 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3294_ (
  .in1({ S248, S5926 }),
  .out1({ S2728 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3295_ (
  .in1({ S249, new_datapath_addsubunit_in1_5 }),
  .out1({ S2729 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3296_ (
  .in1({ S2728, S2598 }),
  .out1({ S2730 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3297_ (
  .in1({ S2729, S2599 }),
  .out1({ S2731 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3298_ (
  .in1({ S240, S5926 }),
  .out1({ S2732 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3299_ (
  .in1({ S241, new_datapath_addsubunit_in1_5 }),
  .out1({ S2733 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3300_ (
  .in1({ S2729, S2599 }),
  .out1({ S2735 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3301_ (
  .in1({ S2728, S2598 }),
  .out1({ S2736 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3302_ (
  .in1({ S2735, S2730 }),
  .out1({ S2737 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3303_ (
  .in1({ S2736, S2731 }),
  .out1({ S2738 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3304_ (
  .in1({ S2738, S2727 }),
  .out1({ S2739 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3305_ (
  .in1({ S2737, S2726 }),
  .out1({ S2740 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3306_ (
  .in1({ S2737, S2726 }),
  .out1({ S2741 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3307_ (
  .in1({ S2738, S2727 }),
  .out1({ S2742 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3308_ (
  .in1({ S2741, S2739 }),
  .out1({ S2743 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3309_ (
  .in1({ S2742, S2740 }),
  .out1({ S2744 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3310_ (
  .in1({ S2623, S2619 }),
  .out1({ S2746 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3311_ (
  .in1({ S2624, S2620 }),
  .out1({ S2747 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3312_ (
  .in1({ S256, S5916 }),
  .out1({ S2748 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3313_ (
  .in1({ S257, new_datapath_addsubunit_in1_6 }),
  .out1({ S2749 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3314_ (
  .in1({ S271, new_datapath_addsubunit_in1_8 }),
  .out1({ S2750 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3315_ (
  .in1({ S2750, S2618 }),
  .out1({ S2751 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3316_ (
  .in1({ S2751 }),
  .out1({ S2752 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3317_ (
  .in1({ S264, S3325 }),
  .out1({ S2753 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3318_ (
  .in1({ S265, new_datapath_addsubunit_in1_8 }),
  .out1({ S2754 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3319_ (
  .in1({ S2754, S887 }),
  .out1({ S2755 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3320_ (
  .in1({ S2753, S886 }),
  .out1({ S2757 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3321_ (
  .in1({ S2755, S2752 }),
  .out1({ S2758 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3322_ (
  .in1({ S2757, S2751 }),
  .out1({ S2759 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3323_ (
  .in1({ S2759, S2749 }),
  .out1({ S2760 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3324_ (
  .in1({ S2758, S2748 }),
  .out1({ S2761 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3325_ (
  .in1({ S2758, S2748 }),
  .out1({ S2762 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3326_ (
  .in1({ S2759, S2749 }),
  .out1({ S2763 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3327_ (
  .in1({ S2762, S2760 }),
  .out1({ S2764 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3328_ (
  .in1({ S2763, S2761 }),
  .out1({ S2765 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3329_ (
  .in1({ S2765, S2746 }),
  .out1({ S2766 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3330_ (
  .in1({ S2764, S2747 }),
  .out1({ S2768 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3331_ (
  .in1({ S2764, S2747 }),
  .out1({ S2769 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3332_ (
  .in1({ S2765, S2746 }),
  .out1({ S2770 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3333_ (
  .in1({ S2769, S2766 }),
  .out1({ S2771 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3334_ (
  .in1({ S2770, S2768 }),
  .out1({ S2772 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3335_ (
  .in1({ S2772, S2744 }),
  .out1({ S2773 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3336_ (
  .in1({ S2771, S2743 }),
  .out1({ S2774 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3337_ (
  .in1({ S2771, S2743 }),
  .out1({ S2775 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3338_ (
  .in1({ S2772, S2744 }),
  .out1({ S2776 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3339_ (
  .in1({ S2775, S2773 }),
  .out1({ S2777 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3340_ (
  .in1({ S2776, S2774 }),
  .out1({ S2779 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3341_ (
  .in1({ S2779, S2724 }),
  .out1({ S2780 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3342_ (
  .in1({ S2777, S2725 }),
  .out1({ S2781 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3343_ (
  .in1({ S2777, S2725 }),
  .out1({ S2782 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3344_ (
  .in1({ S2779, S2724 }),
  .out1({ S2783 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3345_ (
  .in1({ S2782, S2780 }),
  .out1({ S2784 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3346_ (
  .in1({ S2783, S2781 }),
  .out1({ S2785 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3347_ (
  .in1({ S2785, S2722 }),
  .out1({ S2786 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3348_ (
  .in1({ S2784, S2721 }),
  .out1({ S2787 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3349_ (
  .in1({ S2784, S2721 }),
  .out1({ S2788 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3350_ (
  .in1({ S2785, S2722 }),
  .out1({ S2790 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3351_ (
  .in1({ S2788, S2786 }),
  .out1({ S2791 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3352_ (
  .in1({ S2790, S2787 }),
  .out1({ S2792 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3353_ (
  .in1({ S2792, S2686 }),
  .out1({ S2793 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3354_ (
  .in1({ S2791, S2687 }),
  .out1({ S2794 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3355_ (
  .in1({ S2791, S2687 }),
  .out1({ S2795 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3356_ (
  .in1({ S2792, S2686 }),
  .out1({ S2796 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3357_ (
  .in1({ S2795, S2793 }),
  .out1({ S2797 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3358_ (
  .in1({ S2796, S2794 }),
  .out1({ S2798 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3359_ (
  .in1({ S2798, S2586 }),
  .out1({ S2799 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3360_ (
  .in1({ S2797, S2585 }),
  .out1({ S2801 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3361_ (
  .in1({ S2797, S2585 }),
  .out1({ S2802 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3362_ (
  .in1({ S2798, S2586 }),
  .out1({ S2803 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3363_ (
  .in1({ S2802, S2799 }),
  .out1({ S2804 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3364_ (
  .in1({ S2803, S2801 }),
  .out1({ S2805 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3365_ (
  .in1({ S2805, S2684 }),
  .out1({ S2806 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3366_ (
  .in1({ S2805, S2684 }),
  .out1({ S2807 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3367_ (
  .in1({ S2804, S2685 }),
  .out1({ S2808 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3368_ (
  .in1({ S2808, S2806 }),
  .out1({ S2809 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3369_ (
  .in1({ S2809 }),
  .out1({ S2810 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3370_ (
  .in1({ S2810, S2668 }),
  .out1({ S2812 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3371_ (
  .in1({ S2812 }),
  .out1({ S2813 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3372_ (
  .in1({ S2809, S2667 }),
  .out1({ S2814 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3373_ (
  .in1({ S2814, S2812 }),
  .out1({ S2815 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3374_ (
  .in1({ S2815, S2677 }),
  .out1({ S2816 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3375_ (
  .in1({ S2816 }),
  .out1({ S2817 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3376_ (
  .in1({ S2815, S2677 }),
  .out1({ S2818 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3377_ (
  .in1({ S2818, S2817 }),
  .out1({ S2819 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3378_ (
  .in1({ S2819, S2673 }),
  .out1({ S2820 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3379_ (
  .in1({ S2819, S2673 }),
  .out1({ S2821 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3380_ (
  .in1({ S2821, S5579 }),
  .out1({ S2823 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3381_ (
  .in1({ S2823, S2820 }),
  .out1({ S2824 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3382_ (
  .in1({ S2824, S2682 }),
  .out1({ S2825 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3383_ (
  .in1({ S2825, S2683 }),
  .out1({ S28 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3384_ (
  .in1({ S664, S5547 }),
  .out1({ S2826 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3385_ (
  .in1({ S5611, new_datapath_multdivunit_outmdu1_9 }),
  .out1({ S2827 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3386_ (
  .in1({ S2820, S2816 }),
  .out1({ S2828 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3387_ (
  .in1({ S2799, S2793 }),
  .out1({ S2829 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3388_ (
  .in1({ S2801, S2794 }),
  .out1({ S2830 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3389_ (
  .in1({ S5975, S3467 }),
  .out1({ S2831 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3390_ (
  .in1({ new_datapath_addsubunit_in1_0, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S2833 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3391_ (
  .in1({ S2717, S2710 }),
  .out1({ S2834 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3392_ (
  .in1({ S2718, S2711 }),
  .out1({ S2835 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3393_ (
  .in1({ S2834, S2833 }),
  .out1({ S2836 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3394_ (
  .in1({ S2835, S2831 }),
  .out1({ S2837 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3395_ (
  .in1({ S2835, S2831 }),
  .out1({ S2838 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3396_ (
  .in1({ S2834, S2833 }),
  .out1({ S2839 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3397_ (
  .in1({ S2838, S2836 }),
  .out1({ S2840 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3398_ (
  .in1({ S2839, S2837 }),
  .out1({ S2841 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3399_ (
  .in1({ S2786, S2780 }),
  .out1({ S2842 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3400_ (
  .in1({ S2787, S2781 }),
  .out1({ S2844 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3401_ (
  .in1({ S2702, S2697 }),
  .out1({ S2845 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3402_ (
  .in1({ S2703, S2698 }),
  .out1({ S2846 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3403_ (
  .in1({ S5966, S3478 }),
  .out1({ S2847 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3404_ (
  .in1({ new_datapath_addsubunit_in1_1, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S2848 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3405_ (
  .in1({ S202, S5947 }),
  .out1({ S2849 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3406_ (
  .in1({ S203, new_datapath_addsubunit_in1_3 }),
  .out1({ S2850 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3407_ (
  .in1({ S2849, S2695 }),
  .out1({ S2851 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3408_ (
  .in1({ S2850, S2696 }),
  .out1({ S2852 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3409_ (
  .in1({ S228, S5947 }),
  .out1({ S2853 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3410_ (
  .in1({ S229, new_datapath_addsubunit_in1_3 }),
  .out1({ S2855 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3411_ (
  .in1({ S2850, S2696 }),
  .out1({ S2856 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3412_ (
  .in1({ S2849, S2695 }),
  .out1({ S2857 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3413_ (
  .in1({ S2856, S2851 }),
  .out1({ S2858 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3414_ (
  .in1({ S2857, S2852 }),
  .out1({ S2859 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3415_ (
  .in1({ S2859, S2848 }),
  .out1({ S2860 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3416_ (
  .in1({ S2858, S2847 }),
  .out1({ S2861 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3417_ (
  .in1({ S2858, S2847 }),
  .out1({ S2862 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3418_ (
  .in1({ S2859, S2848 }),
  .out1({ S2863 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3419_ (
  .in1({ S2862, S2860 }),
  .out1({ S2864 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3420_ (
  .in1({ S2863, S2861 }),
  .out1({ S2866 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3421_ (
  .in1({ S2739, S2735 }),
  .out1({ S2867 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3422_ (
  .in1({ S2740, S2736 }),
  .out1({ S2868 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3423_ (
  .in1({ S2867, S2866 }),
  .out1({ S2869 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3424_ (
  .in1({ S2868, S2864 }),
  .out1({ S2870 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3425_ (
  .in1({ S2868, S2864 }),
  .out1({ S2871 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3426_ (
  .in1({ S2867, S2866 }),
  .out1({ S2872 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3427_ (
  .in1({ S2871, S2869 }),
  .out1({ S2873 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3428_ (
  .in1({ S2872, S2870 }),
  .out1({ S2874 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3429_ (
  .in1({ S2873, S2846 }),
  .out1({ S2875 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3430_ (
  .in1({ S2874, S2845 }),
  .out1({ S2877 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3431_ (
  .in1({ S2874, S2845 }),
  .out1({ S2878 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3432_ (
  .in1({ S2873, S2846 }),
  .out1({ S2879 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3433_ (
  .in1({ S2878, S2875 }),
  .out1({ S2880 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3434_ (
  .in1({ S2879, S2877 }),
  .out1({ S2881 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3435_ (
  .in1({ S2773, S2766 }),
  .out1({ S2882 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3436_ (
  .in1({ S2774, S2768 }),
  .out1({ S2883 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3437_ (
  .in1({ S208, S5936 }),
  .out1({ S2884 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3438_ (
  .in1({ S209, new_datapath_addsubunit_in1_4 }),
  .out1({ S2885 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3439_ (
  .in1({ S248, S5916 }),
  .out1({ S2886 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3440_ (
  .in1({ S249, new_datapath_addsubunit_in1_6 }),
  .out1({ S2888 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3441_ (
  .in1({ S2886, S2732 }),
  .out1({ S2889 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3442_ (
  .in1({ S2888, S2733 }),
  .out1({ S2890 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3443_ (
  .in1({ S240, S5916 }),
  .out1({ S2891 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3444_ (
  .in1({ S241, new_datapath_addsubunit_in1_6 }),
  .out1({ S2892 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3445_ (
  .in1({ S2888, S2733 }),
  .out1({ S2893 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3446_ (
  .in1({ S2886, S2732 }),
  .out1({ S2894 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3447_ (
  .in1({ S2893, S2889 }),
  .out1({ S2895 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3448_ (
  .in1({ S2894, S2890 }),
  .out1({ S2896 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3449_ (
  .in1({ S2896, S2885 }),
  .out1({ S2897 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3450_ (
  .in1({ S2895, S2884 }),
  .out1({ S2899 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3451_ (
  .in1({ S2895, S2884 }),
  .out1({ S2900 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3452_ (
  .in1({ S2896, S2885 }),
  .out1({ S2901 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3453_ (
  .in1({ S2900, S2897 }),
  .out1({ S2902 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3454_ (
  .in1({ S2901, S2899 }),
  .out1({ S2903 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3455_ (
  .in1({ S2760, S2755 }),
  .out1({ S2904 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3456_ (
  .in1({ S2761, S2757 }),
  .out1({ S2905 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3457_ (
  .in1({ S256, S5907 }),
  .out1({ S2906 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3458_ (
  .in1({ S257, new_datapath_addsubunit_in1_7 }),
  .out1({ S2907 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3459_ (
  .in1({ S2753, S736 }),
  .out1({ S2908 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3460_ (
  .in1({ S2754, S737 }),
  .out1({ S2910 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3461_ (
  .in1({ S265, new_datapath_addsubunit_in1_9 }),
  .out1({ S2911 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3462_ (
  .in1({ S2754, S737 }),
  .out1({ S2912 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3463_ (
  .in1({ S2753, S736 }),
  .out1({ S2913 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3464_ (
  .in1({ S2912, S2908 }),
  .out1({ S2914 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3465_ (
  .in1({ S2913, S2910 }),
  .out1({ S2915 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3466_ (
  .in1({ S2915, S2907 }),
  .out1({ S2916 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3467_ (
  .in1({ S2914, S2906 }),
  .out1({ S2917 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3468_ (
  .in1({ S2914, S2906 }),
  .out1({ S2918 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3469_ (
  .in1({ S2915, S2907 }),
  .out1({ S2919 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3470_ (
  .in1({ S2918, S2916 }),
  .out1({ S2921 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3471_ (
  .in1({ S2919, S2917 }),
  .out1({ S2922 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3472_ (
  .in1({ S2922, S2904 }),
  .out1({ S2923 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3473_ (
  .in1({ S2921, S2905 }),
  .out1({ S2924 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3474_ (
  .in1({ S2921, S2905 }),
  .out1({ S2925 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3475_ (
  .in1({ S2922, S2904 }),
  .out1({ S2926 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3476_ (
  .in1({ S2925, S2923 }),
  .out1({ S2927 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3477_ (
  .in1({ S2926, S2924 }),
  .out1({ S2928 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3478_ (
  .in1({ S2928, S2903 }),
  .out1({ S2929 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3479_ (
  .in1({ S2927, S2902 }),
  .out1({ S2930 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3480_ (
  .in1({ S2927, S2902 }),
  .out1({ S2932 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3481_ (
  .in1({ S2928, S2903 }),
  .out1({ S2933 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3482_ (
  .in1({ S2932, S2929 }),
  .out1({ S2934 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3483_ (
  .in1({ S2933, S2930 }),
  .out1({ S2935 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3484_ (
  .in1({ S2935, S2882 }),
  .out1({ S2936 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3485_ (
  .in1({ S2934, S2883 }),
  .out1({ S2937 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3486_ (
  .in1({ S2934, S2883 }),
  .out1({ S2938 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3487_ (
  .in1({ S2935, S2882 }),
  .out1({ S2939 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3488_ (
  .in1({ S2938, S2936 }),
  .out1({ S2940 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3489_ (
  .in1({ S2939, S2937 }),
  .out1({ S2941 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3490_ (
  .in1({ S2941, S2881 }),
  .out1({ S2943 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3491_ (
  .in1({ S2940, S2880 }),
  .out1({ S2944 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3492_ (
  .in1({ S2940, S2880 }),
  .out1({ S2945 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3493_ (
  .in1({ S2941, S2881 }),
  .out1({ S2946 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3494_ (
  .in1({ S2945, S2943 }),
  .out1({ S2947 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3495_ (
  .in1({ S2946, S2944 }),
  .out1({ S2948 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3496_ (
  .in1({ S2948, S2842 }),
  .out1({ S2949 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3497_ (
  .in1({ S2947, S2844 }),
  .out1({ S2950 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3498_ (
  .in1({ S2947, S2844 }),
  .out1({ S2951 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3499_ (
  .in1({ S2948, S2842 }),
  .out1({ S2952 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3500_ (
  .in1({ S2951, S2949 }),
  .out1({ S2954 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3501_ (
  .in1({ S2952, S2950 }),
  .out1({ S2955 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3502_ (
  .in1({ S2955, S2841 }),
  .out1({ S2956 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3503_ (
  .in1({ S2954, S2840 }),
  .out1({ S2957 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3504_ (
  .in1({ S2954, S2840 }),
  .out1({ S2958 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3505_ (
  .in1({ S2955, S2841 }),
  .out1({ S2959 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3506_ (
  .in1({ S2958, S2956 }),
  .out1({ S2960 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3507_ (
  .in1({ S2959, S2957 }),
  .out1({ S2961 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3508_ (
  .in1({ S2960, S2830 }),
  .out1({ S2962 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3509_ (
  .in1({ S2961, S2829 }),
  .out1({ S2963 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3510_ (
  .in1({ S2961, S2829 }),
  .out1({ S2965 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3511_ (
  .in1({ S2965 }),
  .out1({ S2966 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3512_ (
  .in1({ S2965, S2962 }),
  .out1({ S2967 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3513_ (
  .in1({ S2966, S2963 }),
  .out1({ S2968 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3514_ (
  .in1({ S2968, S2808 }),
  .out1({ S2969 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3515_ (
  .in1({ S2967, S2807 }),
  .out1({ S2970 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3516_ (
  .in1({ S2967, S2807 }),
  .out1({ S2971 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3517_ (
  .in1({ S2968, S2808 }),
  .out1({ S2972 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3518_ (
  .in1({ S2971, S2969 }),
  .out1({ S2973 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3519_ (
  .in1({ S2972, S2970 }),
  .out1({ S2974 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3520_ (
  .in1({ S2973, S2813 }),
  .out1({ S2976 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3521_ (
  .in1({ S2974, S2812 }),
  .out1({ S2977 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3522_ (
  .in1({ S2977, S2976 }),
  .out1({ S2978 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3523_ (
  .in1({ S2978, S2828 }),
  .out1({ S2979 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3524_ (
  .in1({ S2979 }),
  .out1({ S2980 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3525_ (
  .in1({ S2978, S2828 }),
  .out1({ S2981 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3526_ (
  .in1({ S2981, S5579 }),
  .out1({ S2982 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3527_ (
  .in1({ S2982, S2979 }),
  .out1({ S2983 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3528_ (
  .in1({ S2983, S2826 }),
  .out1({ S2984 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3529_ (
  .in1({ S2984, S2827 }),
  .out1({ S29 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3530_ (
  .in1({ S557, S5547 }),
  .out1({ S2986 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3531_ (
  .in1({ S5611, new_datapath_multdivunit_outmdu1_10 }),
  .out1({ S2987 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3532_ (
  .in1({ S2980, S2976 }),
  .out1({ S2988 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3533_ (
  .in1({ S2956, S2949 }),
  .out1({ S2989 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3534_ (
  .in1({ S2957, S2950 }),
  .out1({ S2990 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3535_ (
  .in1({ new_datapath_addsubunit_in1_0, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S2991 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3536_ (
  .in1({ new_datapath_addsubunit_in1_1, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S2992 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3537_ (
  .in1({ S2992, S2991 }),
  .out1({ S2993 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3538_ (
  .in1({ S2993 }),
  .out1({ S2994 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3539_ (
  .in1({ S5966, S3456 }),
  .out1({ S2995 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3540_ (
  .in1({ new_datapath_addsubunit_in1_1, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S2997 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3541_ (
  .in1({ S2997, S2833 }),
  .out1({ S2998 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3542_ (
  .in1({ S2995, S2831 }),
  .out1({ S2999 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3543_ (
  .in1({ S2998, S2994 }),
  .out1({ S3000 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3544_ (
  .in1({ S2999, S2993 }),
  .out1({ S3001 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3545_ (
  .in1({ S2878, S2869 }),
  .out1({ S3002 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3546_ (
  .in1({ S2879, S2870 }),
  .out1({ S3003 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3547_ (
  .in1({ S3003, S3000 }),
  .out1({ S3004 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3548_ (
  .in1({ S3002, S3001 }),
  .out1({ S3005 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3549_ (
  .in1({ S3002, S3001 }),
  .out1({ S3006 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3550_ (
  .in1({ S3003, S3000 }),
  .out1({ S3008 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3551_ (
  .in1({ S3006, S3004 }),
  .out1({ S3009 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3552_ (
  .in1({ S3008, S3005 }),
  .out1({ S3010 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3553_ (
  .in1({ S2943, S2936 }),
  .out1({ S3011 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3554_ (
  .in1({ S2944, S2937 }),
  .out1({ S3012 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3555_ (
  .in1({ S2860, S2856 }),
  .out1({ S3013 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3556_ (
  .in1({ S2861, S2857 }),
  .out1({ S3014 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3557_ (
  .in1({ S5957, S3478 }),
  .out1({ S3015 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3558_ (
  .in1({ new_datapath_addsubunit_in1_2, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S3016 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3559_ (
  .in1({ S202, S5936 }),
  .out1({ S3017 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3560_ (
  .in1({ S203, new_datapath_addsubunit_in1_4 }),
  .out1({ S3019 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3561_ (
  .in1({ S3017, S2853 }),
  .out1({ S3020 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3562_ (
  .in1({ S3019, S2855 }),
  .out1({ S3021 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3563_ (
  .in1({ S228, S5936 }),
  .out1({ S3022 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3564_ (
  .in1({ S229, new_datapath_addsubunit_in1_4 }),
  .out1({ S3023 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3565_ (
  .in1({ S3019, S2855 }),
  .out1({ S3024 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3566_ (
  .in1({ S3017, S2853 }),
  .out1({ S3025 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3567_ (
  .in1({ S3024, S3020 }),
  .out1({ S3026 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3568_ (
  .in1({ S3025, S3021 }),
  .out1({ S3027 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3569_ (
  .in1({ S3027, S3016 }),
  .out1({ S3028 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3570_ (
  .in1({ S3026, S3015 }),
  .out1({ S3030 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3571_ (
  .in1({ S3026, S3015 }),
  .out1({ S3031 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3572_ (
  .in1({ S3027, S3016 }),
  .out1({ S3032 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3573_ (
  .in1({ S3031, S3028 }),
  .out1({ S3033 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3574_ (
  .in1({ S3032, S3030 }),
  .out1({ S3034 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3575_ (
  .in1({ S2897, S2893 }),
  .out1({ S3035 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3576_ (
  .in1({ S2899, S2894 }),
  .out1({ S3036 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3577_ (
  .in1({ S3035, S3034 }),
  .out1({ S3037 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3578_ (
  .in1({ S3036, S3033 }),
  .out1({ S3038 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3579_ (
  .in1({ S3036, S3033 }),
  .out1({ S3039 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3580_ (
  .in1({ S3035, S3034 }),
  .out1({ S3041 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3581_ (
  .in1({ S3039, S3037 }),
  .out1({ S3042 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3582_ (
  .in1({ S3041, S3038 }),
  .out1({ S3043 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3583_ (
  .in1({ S3042, S3014 }),
  .out1({ S3044 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3584_ (
  .in1({ S3043, S3013 }),
  .out1({ S3045 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3585_ (
  .in1({ S3043, S3013 }),
  .out1({ S3046 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3586_ (
  .in1({ S3042, S3014 }),
  .out1({ S3047 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3587_ (
  .in1({ S3046, S3044 }),
  .out1({ S3048 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3588_ (
  .in1({ S3047, S3045 }),
  .out1({ S3049 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3589_ (
  .in1({ S2929, S2923 }),
  .out1({ S3050 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3590_ (
  .in1({ S2930, S2924 }),
  .out1({ S3052 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3591_ (
  .in1({ S208, S5926 }),
  .out1({ S3053 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3592_ (
  .in1({ S209, new_datapath_addsubunit_in1_5 }),
  .out1({ S3054 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3593_ (
  .in1({ S248, S5907 }),
  .out1({ S3055 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3594_ (
  .in1({ S249, new_datapath_addsubunit_in1_7 }),
  .out1({ S3056 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3595_ (
  .in1({ S3055, S2891 }),
  .out1({ S3057 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3596_ (
  .in1({ S3056, S2892 }),
  .out1({ S3058 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3597_ (
  .in1({ S240, S5907 }),
  .out1({ S3059 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3598_ (
  .in1({ S241, new_datapath_addsubunit_in1_7 }),
  .out1({ S3060 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3599_ (
  .in1({ S3056, S2892 }),
  .out1({ S3061 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3600_ (
  .in1({ S3055, S2891 }),
  .out1({ S3063 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3601_ (
  .in1({ S3061, S3057 }),
  .out1({ S3064 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3602_ (
  .in1({ S3063, S3058 }),
  .out1({ S3065 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3603_ (
  .in1({ S3065, S3054 }),
  .out1({ S3066 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3604_ (
  .in1({ S3064, S3053 }),
  .out1({ S3067 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3605_ (
  .in1({ S3064, S3053 }),
  .out1({ S3068 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3606_ (
  .in1({ S3065, S3054 }),
  .out1({ S3069 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3607_ (
  .in1({ S3068, S3066 }),
  .out1({ S3070 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3608_ (
  .in1({ S3069, S3067 }),
  .out1({ S3071 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3609_ (
  .in1({ S2916, S2912 }),
  .out1({ S3072 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3610_ (
  .in1({ S2917, S2913 }),
  .out1({ S3074 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3611_ (
  .in1({ S257, new_datapath_addsubunit_in1_8 }),
  .out1({ S3075 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3612_ (
  .in1({ S3075 }),
  .out1({ S3076 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3613_ (
  .in1({ S271, new_datapath_addsubunit_in1_10 }),
  .out1({ S3077 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3614_ (
  .in1({ S3077, S2911 }),
  .out1({ S3078 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3615_ (
  .in1({ S264, S3346 }),
  .out1({ S3079 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3616_ (
  .in1({ S265, new_datapath_addsubunit_in1_10 }),
  .out1({ S3080 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3617_ (
  .in1({ S3080, S737 }),
  .out1({ S3081 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3618_ (
  .in1({ S3079, S736 }),
  .out1({ S3082 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3619_ (
  .in1({ S3082, S3078 }),
  .out1({ S3083 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3620_ (
  .in1({ S3083 }),
  .out1({ S3085 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3621_ (
  .in1({ S3083, S3075 }),
  .out1({ S3086 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3622_ (
  .in1({ S3085, S3076 }),
  .out1({ S3087 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3623_ (
  .in1({ S3083, S3075 }),
  .out1({ S3088 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3624_ (
  .in1({ S3088 }),
  .out1({ S3089 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3625_ (
  .in1({ S3089, S3086 }),
  .out1({ S3090 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3626_ (
  .in1({ S3088, S3087 }),
  .out1({ S3091 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3627_ (
  .in1({ S3091, S3072 }),
  .out1({ S3092 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3628_ (
  .in1({ S3090, S3074 }),
  .out1({ S3093 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3629_ (
  .in1({ S3090, S3074 }),
  .out1({ S3094 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3630_ (
  .in1({ S3091, S3072 }),
  .out1({ S3096 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3631_ (
  .in1({ S3094, S3092 }),
  .out1({ S3097 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3632_ (
  .in1({ S3096, S3093 }),
  .out1({ S3098 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3633_ (
  .in1({ S3098, S3071 }),
  .out1({ S3099 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3634_ (
  .in1({ S3097, S3070 }),
  .out1({ S3100 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3635_ (
  .in1({ S3097, S3070 }),
  .out1({ S3101 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3636_ (
  .in1({ S3098, S3071 }),
  .out1({ S3102 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3637_ (
  .in1({ S3101, S3099 }),
  .out1({ S3103 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3638_ (
  .in1({ S3102, S3100 }),
  .out1({ S3104 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3639_ (
  .in1({ S3104, S3050 }),
  .out1({ S3105 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3640_ (
  .in1({ S3103, S3052 }),
  .out1({ S3107 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3641_ (
  .in1({ S3103, S3052 }),
  .out1({ S3108 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3642_ (
  .in1({ S3104, S3050 }),
  .out1({ S3109 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3643_ (
  .in1({ S3108, S3105 }),
  .out1({ S3110 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3644_ (
  .in1({ S3109, S3107 }),
  .out1({ S3111 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3645_ (
  .in1({ S3111, S3049 }),
  .out1({ S3112 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3646_ (
  .in1({ S3110, S3048 }),
  .out1({ S3113 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3647_ (
  .in1({ S3110, S3048 }),
  .out1({ S3114 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3648_ (
  .in1({ S3111, S3049 }),
  .out1({ S3115 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3649_ (
  .in1({ S3114, S3112 }),
  .out1({ S3116 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3650_ (
  .in1({ S3115, S3113 }),
  .out1({ S3118 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3651_ (
  .in1({ S3118, S3011 }),
  .out1({ S3119 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3652_ (
  .in1({ S3116, S3012 }),
  .out1({ S3120 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3653_ (
  .in1({ S3116, S3012 }),
  .out1({ S3121 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3654_ (
  .in1({ S3118, S3011 }),
  .out1({ S3122 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3655_ (
  .in1({ S3121, S3119 }),
  .out1({ S3123 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3656_ (
  .in1({ S3122, S3120 }),
  .out1({ S3124 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3657_ (
  .in1({ S3124, S3010 }),
  .out1({ S3125 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3658_ (
  .in1({ S3123, S3009 }),
  .out1({ S3126 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3659_ (
  .in1({ S3123, S3009 }),
  .out1({ S3127 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3660_ (
  .in1({ S3124, S3010 }),
  .out1({ S3129 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3661_ (
  .in1({ S3127, S3125 }),
  .out1({ S3130 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3662_ (
  .in1({ S3129, S3126 }),
  .out1({ S3131 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3663_ (
  .in1({ S3131, S2989 }),
  .out1({ S3132 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3664_ (
  .in1({ S3130, S2990 }),
  .out1({ S3133 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3665_ (
  .in1({ S3130, S2990 }),
  .out1({ S3134 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3666_ (
  .in1({ S3131, S2989 }),
  .out1({ S3135 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3667_ (
  .in1({ S3134, S3132 }),
  .out1({ S3136 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3668_ (
  .in1({ S3135, S3133 }),
  .out1({ S3137 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3669_ (
  .in1({ S3137, S2837 }),
  .out1({ S3138 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3670_ (
  .in1({ S3136, S2836 }),
  .out1({ S3140 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3671_ (
  .in1({ S3140, S3138 }),
  .out1({ S3141 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3672_ (
  .in1({ S3141, S2965 }),
  .out1({ S3142 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3673_ (
  .in1({ S3142 }),
  .out1({ S3143 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3674_ (
  .in1({ S3141, S2965 }),
  .out1({ S3144 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3675_ (
  .in1({ S3144 }),
  .out1({ S3145 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3676_ (
  .in1({ S3144, S3143 }),
  .out1({ S3146 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3677_ (
  .in1({ S3145, S3142 }),
  .out1({ S3147 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3678_ (
  .in1({ S3147, S2970 }),
  .out1({ S3148 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3679_ (
  .in1({ S3146, S2969 }),
  .out1({ S3149 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3680_ (
  .in1({ S3149, S3148 }),
  .out1({ S3151 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3681_ (
  .in1({ S3151, S2988 }),
  .out1({ S3152 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3682_ (
  .in1({ S3152 }),
  .out1({ S3153 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3683_ (
  .in1({ S3151, S2988 }),
  .out1({ S3154 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3684_ (
  .in1({ S3152, S5579 }),
  .out1({ S3155 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3685_ (
  .in1({ S3155, S3154 }),
  .out1({ S3156 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3686_ (
  .in1({ S3156, S2986 }),
  .out1({ S3157 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3687_ (
  .in1({ S3157, S2987 }),
  .out1({ S30 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3688_ (
  .in1({ S461, S5547 }),
  .out1({ S3158 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3689_ (
  .in1({ S5611, new_datapath_multdivunit_outmdu1_11 }),
  .out1({ S3159 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3690_ (
  .in1({ S3153, S3148 }),
  .out1({ S3161 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3691_ (
  .in1({ S3138, S3132 }),
  .out1({ S3162 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3692_ (
  .in1({ S3162 }),
  .out1({ S3163 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3693_ (
  .in1({ S3125, S3119 }),
  .out1({ S3164 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3694_ (
  .in1({ S3126, S3120 }),
  .out1({ S3165 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3695_ (
  .in1({ new_datapath_addsubunit_in1_0, new_datapath_multdivunit_1697_B_11 }),
  .out1({ S3166 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3696_ (
  .in1({ S3166 }),
  .out1({ S3167 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3697_ (
  .in1({ S5957, S3467 }),
  .out1({ S3168 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3698_ (
  .in1({ new_datapath_addsubunit_in1_2, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S3169 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3699_ (
  .in1({ S3169, S2997 }),
  .out1({ S3170 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3700_ (
  .in1({ new_datapath_addsubunit_in1_2, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S3172 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3701_ (
  .in1({ S3169, S2997 }),
  .out1({ S3173 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3702_ (
  .in1({ S3168, S2995 }),
  .out1({ S3174 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3703_ (
  .in1({ S3174, S3170 }),
  .out1({ S3175 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3704_ (
  .in1({ S3175 }),
  .out1({ S3176 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3705_ (
  .in1({ S3175, S3166 }),
  .out1({ S3177 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3706_ (
  .in1({ S3176, S3167 }),
  .out1({ S3178 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3707_ (
  .in1({ S3175, S3166 }),
  .out1({ S3179 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3708_ (
  .in1({ S3179 }),
  .out1({ S3180 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3709_ (
  .in1({ S3180, S3177 }),
  .out1({ S3181 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3710_ (
  .in1({ S3179, S3178 }),
  .out1({ S3183 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3711_ (
  .in1({ S3183, S2999 }),
  .out1({ S3184 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3712_ (
  .in1({ S3181, S2998 }),
  .out1({ S3185 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3713_ (
  .in1({ S3181, S2998 }),
  .out1({ S3186 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3714_ (
  .in1({ S3183, S2999 }),
  .out1({ S3187 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3715_ (
  .in1({ S3186, S3184 }),
  .out1({ S3188 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3716_ (
  .in1({ S3187, S3185 }),
  .out1({ S3189 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3717_ (
  .in1({ S3046, S3037 }),
  .out1({ S3190 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3718_ (
  .in1({ S3047, S3038 }),
  .out1({ S3191 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3719_ (
  .in1({ S3191, S3188 }),
  .out1({ S3192 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3720_ (
  .in1({ S3190, S3189 }),
  .out1({ S3194 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3721_ (
  .in1({ S3190, S3189 }),
  .out1({ S3195 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3722_ (
  .in1({ S3191, S3188 }),
  .out1({ S3196 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3723_ (
  .in1({ S3195, S3192 }),
  .out1({ S3197 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3724_ (
  .in1({ S3196, S3194 }),
  .out1({ S3198 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3725_ (
  .in1({ S3112, S3105 }),
  .out1({ S3199 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3726_ (
  .in1({ S3113, S3107 }),
  .out1({ S3200 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3727_ (
  .in1({ S3028, S3024 }),
  .out1({ S3201 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3728_ (
  .in1({ S3030, S3025 }),
  .out1({ S3202 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3729_ (
  .in1({ S5947, S3478 }),
  .out1({ S3203 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3730_ (
  .in1({ new_datapath_addsubunit_in1_3, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S3205 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3731_ (
  .in1({ S202, S5926 }),
  .out1({ S3206 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3732_ (
  .in1({ S203, new_datapath_addsubunit_in1_5 }),
  .out1({ S3207 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3733_ (
  .in1({ S3206, S3022 }),
  .out1({ S3208 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3734_ (
  .in1({ S3207, S3023 }),
  .out1({ S3209 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3735_ (
  .in1({ S228, S5926 }),
  .out1({ S3210 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3736_ (
  .in1({ S229, new_datapath_addsubunit_in1_5 }),
  .out1({ S3211 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3737_ (
  .in1({ S3207, S3023 }),
  .out1({ S3212 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3738_ (
  .in1({ S3206, S3022 }),
  .out1({ S3213 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3739_ (
  .in1({ S3212, S3208 }),
  .out1({ S3214 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3740_ (
  .in1({ S3213, S3209 }),
  .out1({ S3216 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3741_ (
  .in1({ S3216, S3205 }),
  .out1({ S3217 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3742_ (
  .in1({ S3214, S3203 }),
  .out1({ S3218 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3743_ (
  .in1({ S3214, S3203 }),
  .out1({ S3219 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3744_ (
  .in1({ S3216, S3205 }),
  .out1({ S3220 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3745_ (
  .in1({ S3219, S3217 }),
  .out1({ S3221 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3746_ (
  .in1({ S3220, S3218 }),
  .out1({ S3222 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3747_ (
  .in1({ S3066, S3061 }),
  .out1({ S3223 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3748_ (
  .in1({ S3067, S3063 }),
  .out1({ S3224 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3749_ (
  .in1({ S3223, S3222 }),
  .out1({ S3225 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3750_ (
  .in1({ S3224, S3221 }),
  .out1({ S3227 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3751_ (
  .in1({ S3224, S3221 }),
  .out1({ S3228 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3752_ (
  .in1({ S3223, S3222 }),
  .out1({ S3229 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3753_ (
  .in1({ S3228, S3225 }),
  .out1({ S3230 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3754_ (
  .in1({ S3229, S3227 }),
  .out1({ S3231 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3755_ (
  .in1({ S3230, S3202 }),
  .out1({ S3232 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3756_ (
  .in1({ S3231, S3201 }),
  .out1({ S3233 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3757_ (
  .in1({ S3231, S3201 }),
  .out1({ S3234 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3758_ (
  .in1({ S3230, S3202 }),
  .out1({ S3235 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3759_ (
  .in1({ S3234, S3232 }),
  .out1({ S3236 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3760_ (
  .in1({ S3235, S3233 }),
  .out1({ S3238 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3761_ (
  .in1({ S3099, S3092 }),
  .out1({ S3239 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3762_ (
  .in1({ S3100, S3093 }),
  .out1({ S3240 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3763_ (
  .in1({ S208, S5916 }),
  .out1({ S3241 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3764_ (
  .in1({ S209, new_datapath_addsubunit_in1_6 }),
  .out1({ S3242 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3765_ (
  .in1({ S248, S3325 }),
  .out1({ S3243 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3766_ (
  .in1({ S249, new_datapath_addsubunit_in1_8 }),
  .out1({ S3244 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3767_ (
  .in1({ S3243, S3059 }),
  .out1({ S3245 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3768_ (
  .in1({ S3244, S3060 }),
  .out1({ S3246 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3769_ (
  .in1({ S241, new_datapath_addsubunit_in1_8 }),
  .out1({ S3247 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3770_ (
  .in1({ S3244, S3060 }),
  .out1({ S3249 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3771_ (
  .in1({ S3243, S3059 }),
  .out1({ S3250 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3772_ (
  .in1({ S3249, S3245 }),
  .out1({ S3251 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3773_ (
  .in1({ S3250, S3246 }),
  .out1({ S3252 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3774_ (
  .in1({ S3252, S3242 }),
  .out1({ S3253 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3775_ (
  .in1({ S3251, S3241 }),
  .out1({ S3254 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3776_ (
  .in1({ S3251, S3241 }),
  .out1({ S3255 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3777_ (
  .in1({ S3252, S3242 }),
  .out1({ S3256 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3778_ (
  .in1({ S3255, S3253 }),
  .out1({ S3257 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3779_ (
  .in1({ S3256, S3254 }),
  .out1({ S3258 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3780_ (
  .in1({ S3086, S3081 }),
  .out1({ S3260 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3781_ (
  .in1({ S3087, S3082 }),
  .out1({ S3261 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3782_ (
  .in1({ S256, S3336 }),
  .out1({ S3262 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3783_ (
  .in1({ S257, new_datapath_addsubunit_in1_9 }),
  .out1({ S3263 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3784_ (
  .in1({ S3079, S511 }),
  .out1({ S3264 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3785_ (
  .in1({ S3080, S512 }),
  .out1({ S3265 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3786_ (
  .in1({ S265, new_datapath_addsubunit_in1_11 }),
  .out1({ S3266 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3787_ (
  .in1({ S3080, S512 }),
  .out1({ S3267 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3788_ (
  .in1({ S3079, S511 }),
  .out1({ S3268 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3789_ (
  .in1({ S3267, S3264 }),
  .out1({ S3269 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3790_ (
  .in1({ S3268, S3265 }),
  .out1({ S3271 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3791_ (
  .in1({ S3271, S3263 }),
  .out1({ S3272 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3792_ (
  .in1({ S3269, S3262 }),
  .out1({ S3273 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3793_ (
  .in1({ S3269, S3262 }),
  .out1({ S3274 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3794_ (
  .in1({ S3271, S3263 }),
  .out1({ S3275 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3795_ (
  .in1({ S3274, S3272 }),
  .out1({ S3276 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3796_ (
  .in1({ S3275, S3273 }),
  .out1({ S3277 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3797_ (
  .in1({ S3277, S3260 }),
  .out1({ S3278 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3798_ (
  .in1({ S3276, S3261 }),
  .out1({ S3279 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3799_ (
  .in1({ S3276, S3261 }),
  .out1({ S3280 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3800_ (
  .in1({ S3277, S3260 }),
  .out1({ S3282 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3801_ (
  .in1({ S3280, S3278 }),
  .out1({ S3283 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3802_ (
  .in1({ S3282, S3279 }),
  .out1({ S3284 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3803_ (
  .in1({ S3284, S3258 }),
  .out1({ S3285 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3804_ (
  .in1({ S3283, S3257 }),
  .out1({ S3286 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3805_ (
  .in1({ S3283, S3257 }),
  .out1({ S3287 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3806_ (
  .in1({ S3284, S3258 }),
  .out1({ S3288 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3807_ (
  .in1({ S3287, S3285 }),
  .out1({ S3289 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3808_ (
  .in1({ S3288, S3286 }),
  .out1({ S3290 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3809_ (
  .in1({ S3290, S3239 }),
  .out1({ S3291 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3810_ (
  .in1({ S3289, S3240 }),
  .out1({ S3293 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3811_ (
  .in1({ S3289, S3240 }),
  .out1({ S3294 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3812_ (
  .in1({ S3290, S3239 }),
  .out1({ S3295 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3813_ (
  .in1({ S3294, S3291 }),
  .out1({ S3296 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3814_ (
  .in1({ S3295, S3293 }),
  .out1({ S3297 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3815_ (
  .in1({ S3297, S3238 }),
  .out1({ S3298 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3816_ (
  .in1({ S3296, S3236 }),
  .out1({ S3299 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3817_ (
  .in1({ S3296, S3236 }),
  .out1({ S3300 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3818_ (
  .in1({ S3297, S3238 }),
  .out1({ S3301 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3819_ (
  .in1({ S3300, S3298 }),
  .out1({ S3302 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3820_ (
  .in1({ S3301, S3299 }),
  .out1({ S3304 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3821_ (
  .in1({ S3304, S3199 }),
  .out1({ S3305 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3822_ (
  .in1({ S3302, S3200 }),
  .out1({ S3306 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3823_ (
  .in1({ S3302, S3200 }),
  .out1({ S3307 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3824_ (
  .in1({ S3304, S3199 }),
  .out1({ S3308 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3825_ (
  .in1({ S3307, S3305 }),
  .out1({ S3309 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3826_ (
  .in1({ S3308, S3306 }),
  .out1({ S3310 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3827_ (
  .in1({ S3310, S3198 }),
  .out1({ S3311 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3828_ (
  .in1({ S3309, S3197 }),
  .out1({ S3312 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3829_ (
  .in1({ S3309, S3197 }),
  .out1({ S3313 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3830_ (
  .in1({ S3310, S3198 }),
  .out1({ S3315 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3831_ (
  .in1({ S3313, S3311 }),
  .out1({ S3316 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3832_ (
  .in1({ S3315, S3312 }),
  .out1({ S3317 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3833_ (
  .in1({ S3317, S3164 }),
  .out1({ S3318 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3834_ (
  .in1({ S3316, S3165 }),
  .out1({ S3319 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3835_ (
  .in1({ S3316, S3165 }),
  .out1({ S3320 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3836_ (
  .in1({ S3317, S3164 }),
  .out1({ S3321 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3837_ (
  .in1({ S3320, S3318 }),
  .out1({ S3322 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3838_ (
  .in1({ S3321, S3319 }),
  .out1({ S3323 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3839_ (
  .in1({ S3323, S3008 }),
  .out1({ S3324 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3840_ (
  .in1({ S3322, S3006 }),
  .out1({ S3326 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3841_ (
  .in1({ S3323, S3008 }),
  .out1({ S3327 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3842_ (
  .in1({ S3327, S3326 }),
  .out1({ S3328 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3843_ (
  .in1({ S3328 }),
  .out1({ S3329 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3844_ (
  .in1({ S3328, S3162 }),
  .out1({ S3330 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3845_ (
  .in1({ S3329, S3163 }),
  .out1({ S3331 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3846_ (
  .in1({ S3331 }),
  .out1({ S3332 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3847_ (
  .in1({ S3331, S3330 }),
  .out1({ S3333 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3848_ (
  .in1({ S3333, S3142 }),
  .out1({ S3334 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3849_ (
  .in1({ S3334 }),
  .out1({ S3335 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3850_ (
  .in1({ S3333, S3142 }),
  .out1({ S3337 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3851_ (
  .in1({ S3337, S3335 }),
  .out1({ S3338 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3852_ (
  .in1({ S3338, S3161 }),
  .out1({ S3339 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3853_ (
  .in1({ S3338, S3161 }),
  .out1({ S3340 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3854_ (
  .in1({ S3340, S5579 }),
  .out1({ S3341 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3855_ (
  .in1({ S3341, S3339 }),
  .out1({ S3342 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3856_ (
  .in1({ S3342, S3158 }),
  .out1({ S3343 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3857_ (
  .in1({ S3343, S3159 }),
  .out1({ S31 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3858_ (
  .in1({ S3339, S3334 }),
  .out1({ S3344 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3859_ (
  .in1({ S3324, S3318 }),
  .out1({ S3345 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3860_ (
  .in1({ S3326, S3319 }),
  .out1({ S3347 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3861_ (
  .in1({ S3311, S3305 }),
  .out1({ S3348 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3862_ (
  .in1({ S3312, S3306 }),
  .out1({ S3349 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3863_ (
  .in1({ S5975, S3434 }),
  .out1({ S3350 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3864_ (
  .in1({ new_datapath_addsubunit_in1_0, new_datapath_multdivunit_1697_B_12 }),
  .out1({ S3351 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3865_ (
  .in1({ S3177, S3173 }),
  .out1({ S3352 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3866_ (
  .in1({ S3178, S3174 }),
  .out1({ S3353 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3867_ (
  .in1({ new_datapath_addsubunit_in1_1, new_datapath_multdivunit_1697_B_11 }),
  .out1({ S3354 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3868_ (
  .in1({ new_datapath_addsubunit_in1_3, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S3355 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3869_ (
  .in1({ S3355, S3172 }),
  .out1({ S3356 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3870_ (
  .in1({ S5947, S3456 }),
  .out1({ S3358 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3871_ (
  .in1({ new_datapath_addsubunit_in1_3, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S3359 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3872_ (
  .in1({ S3355, S3172 }),
  .out1({ S3360 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3873_ (
  .in1({ S3360 }),
  .out1({ S3361 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3874_ (
  .in1({ S3361, S3356 }),
  .out1({ S3362 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3875_ (
  .in1({ S3362, S3354 }),
  .out1({ S3363 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3876_ (
  .in1({ S3363 }),
  .out1({ S3364 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3877_ (
  .in1({ S3362, S3354 }),
  .out1({ S3365 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3878_ (
  .in1({ S3365 }),
  .out1({ S3366 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3879_ (
  .in1({ S3366, S3363 }),
  .out1({ S3367 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3880_ (
  .in1({ S3365, S3364 }),
  .out1({ S3369 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3881_ (
  .in1({ S3369, S3352 }),
  .out1({ S3370 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3882_ (
  .in1({ S3367, S3353 }),
  .out1({ S3371 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3883_ (
  .in1({ S3367, S3353 }),
  .out1({ S3372 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3884_ (
  .in1({ S3369, S3352 }),
  .out1({ S3373 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3885_ (
  .in1({ S3372, S3370 }),
  .out1({ S3374 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3886_ (
  .in1({ S3373, S3371 }),
  .out1({ S3375 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3887_ (
  .in1({ S3375, S3351 }),
  .out1({ S3376 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3888_ (
  .in1({ S3374, S3350 }),
  .out1({ S3377 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3889_ (
  .in1({ S3374, S3350 }),
  .out1({ S3378 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3890_ (
  .in1({ S3375, S3351 }),
  .out1({ S3380 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3891_ (
  .in1({ S3378, S3376 }),
  .out1({ S3381 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3892_ (
  .in1({ S3380, S3377 }),
  .out1({ S3382 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3893_ (
  .in1({ S3234, S3225 }),
  .out1({ S3383 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3894_ (
  .in1({ S3235, S3227 }),
  .out1({ S3384 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3895_ (
  .in1({ S3383, S3382 }),
  .out1({ S3385 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3896_ (
  .in1({ S3384, S3381 }),
  .out1({ S3386 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3897_ (
  .in1({ S3384, S3381 }),
  .out1({ S3387 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3898_ (
  .in1({ S3383, S3382 }),
  .out1({ S3388 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3899_ (
  .in1({ S3387, S3385 }),
  .out1({ S3389 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3900_ (
  .in1({ S3388, S3386 }),
  .out1({ S3391 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3901_ (
  .in1({ S3391, S3185 }),
  .out1({ S3392 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3902_ (
  .in1({ S3389, S3184 }),
  .out1({ S3393 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3903_ (
  .in1({ S3389, S3184 }),
  .out1({ S3394 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3904_ (
  .in1({ S3391, S3185 }),
  .out1({ S3395 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3905_ (
  .in1({ S3394, S3392 }),
  .out1({ S3396 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3906_ (
  .in1({ S3395, S3393 }),
  .out1({ S3397 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3907_ (
  .in1({ S3298, S3291 }),
  .out1({ S3398 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3908_ (
  .in1({ S3299, S3293 }),
  .out1({ S3399 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3909_ (
  .in1({ S3217, S3212 }),
  .out1({ S3400 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3910_ (
  .in1({ S3218, S3213 }),
  .out1({ S3402 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3911_ (
  .in1({ S5936, S3478 }),
  .out1({ S3403 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3912_ (
  .in1({ new_datapath_addsubunit_in1_4, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S3404 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3913_ (
  .in1({ S202, S5916 }),
  .out1({ S3405 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3914_ (
  .in1({ S203, new_datapath_addsubunit_in1_6 }),
  .out1({ S3406 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3915_ (
  .in1({ S3405, S3210 }),
  .out1({ S3407 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3916_ (
  .in1({ S3406, S3211 }),
  .out1({ S3408 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3917_ (
  .in1({ S228, S5916 }),
  .out1({ S3409 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3918_ (
  .in1({ S229, new_datapath_addsubunit_in1_6 }),
  .out1({ S3410 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3919_ (
  .in1({ S3406, S3211 }),
  .out1({ S3411 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3920_ (
  .in1({ S3405, S3210 }),
  .out1({ S3413 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3921_ (
  .in1({ S3411, S3407 }),
  .out1({ S3414 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3922_ (
  .in1({ S3413, S3408 }),
  .out1({ S3415 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3923_ (
  .in1({ S3415, S3404 }),
  .out1({ S3416 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3924_ (
  .in1({ S3414, S3403 }),
  .out1({ S3417 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3925_ (
  .in1({ S3414, S3403 }),
  .out1({ S3418 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3926_ (
  .in1({ S3415, S3404 }),
  .out1({ S3419 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3927_ (
  .in1({ S3418, S3416 }),
  .out1({ S3420 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3928_ (
  .in1({ S3419, S3417 }),
  .out1({ S3421 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3929_ (
  .in1({ S3253, S3249 }),
  .out1({ S3422 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3930_ (
  .in1({ S3254, S3250 }),
  .out1({ S3424 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3931_ (
  .in1({ S3422, S3421 }),
  .out1({ S3425 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3932_ (
  .in1({ S3424, S3420 }),
  .out1({ S3426 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3933_ (
  .in1({ S3424, S3420 }),
  .out1({ S3427 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3934_ (
  .in1({ S3422, S3421 }),
  .out1({ S3428 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3935_ (
  .in1({ S3427, S3425 }),
  .out1({ S3429 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3936_ (
  .in1({ S3428, S3426 }),
  .out1({ S3430 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3937_ (
  .in1({ S3429, S3402 }),
  .out1({ S3431 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3938_ (
  .in1({ S3430, S3400 }),
  .out1({ S3432 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3939_ (
  .in1({ S3430, S3400 }),
  .out1({ S3433 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3940_ (
  .in1({ S3429, S3402 }),
  .out1({ S3435 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3941_ (
  .in1({ S3433, S3431 }),
  .out1({ S3436 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3942_ (
  .in1({ S3435, S3432 }),
  .out1({ S3437 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3943_ (
  .in1({ S3285, S3278 }),
  .out1({ S3438 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3944_ (
  .in1({ S3286, S3279 }),
  .out1({ S3439 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3945_ (
  .in1({ S208, S5907 }),
  .out1({ S3440 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3946_ (
  .in1({ S209, new_datapath_addsubunit_in1_7 }),
  .out1({ S3441 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3947_ (
  .in1({ S249, new_datapath_addsubunit_in1_9 }),
  .out1({ S3442 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3948_ (
  .in1({ S3442, S3247 }),
  .out1({ S3443 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3949_ (
  .in1({ S3443 }),
  .out1({ S3444 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3950_ (
  .in1({ S240, S3336 }),
  .out1({ S3446 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3951_ (
  .in1({ S241, new_datapath_addsubunit_in1_9 }),
  .out1({ S3447 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3952_ (
  .in1({ S3442, S3247 }),
  .out1({ S3448 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3953_ (
  .in1({ S3446, S3243 }),
  .out1({ S3449 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3954_ (
  .in1({ S3448, S3444 }),
  .out1({ S3450 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3955_ (
  .in1({ S3449, S3443 }),
  .out1({ S3451 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3956_ (
  .in1({ S3451, S3441 }),
  .out1({ S3452 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3957_ (
  .in1({ S3450, S3440 }),
  .out1({ S3453 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3958_ (
  .in1({ S3450, S3440 }),
  .out1({ S3454 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3959_ (
  .in1({ S3451, S3441 }),
  .out1({ S3455 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3960_ (
  .in1({ S3454, S3452 }),
  .out1({ S3457 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3961_ (
  .in1({ S3455, S3453 }),
  .out1({ S3458 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3962_ (
  .in1({ S3272, S3267 }),
  .out1({ S3459 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3963_ (
  .in1({ S3273, S3268 }),
  .out1({ S3460 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3964_ (
  .in1({ S257, new_datapath_addsubunit_in1_10 }),
  .out1({ S3461 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3965_ (
  .in1({ S3461 }),
  .out1({ S3462 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3966_ (
  .in1({ S271, new_datapath_addsubunit_in1_12 }),
  .out1({ S3463 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3967_ (
  .in1({ S3463, S3266 }),
  .out1({ S3464 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3968_ (
  .in1({ S264, S3368 }),
  .out1({ S3465 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3969_ (
  .in1({ S265, new_datapath_addsubunit_in1_12 }),
  .out1({ S3466 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3970_ (
  .in1({ S3466, S512 }),
  .out1({ S3468 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3971_ (
  .in1({ S3465, S511 }),
  .out1({ S3469 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3972_ (
  .in1({ S3469, S3464 }),
  .out1({ S3470 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3973_ (
  .in1({ S3470 }),
  .out1({ S3471 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3974_ (
  .in1({ S3470, S3461 }),
  .out1({ S3472 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3975_ (
  .in1({ S3471, S3462 }),
  .out1({ S3473 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3976_ (
  .in1({ S3470, S3461 }),
  .out1({ S3474 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_3977_ (
  .in1({ S3474 }),
  .out1({ S3475 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3978_ (
  .in1({ S3475, S3472 }),
  .out1({ S3476 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3979_ (
  .in1({ S3474, S3473 }),
  .out1({ S3477 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3980_ (
  .in1({ S3477, S3459 }),
  .out1({ S3479 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3981_ (
  .in1({ S3476, S3460 }),
  .out1({ S3480 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3982_ (
  .in1({ S3476, S3460 }),
  .out1({ S3481 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3983_ (
  .in1({ S3477, S3459 }),
  .out1({ S3482 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3984_ (
  .in1({ S3481, S3479 }),
  .out1({ S3483 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3985_ (
  .in1({ S3482, S3480 }),
  .out1({ S3484 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3986_ (
  .in1({ S3484, S3458 }),
  .out1({ S3485 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3987_ (
  .in1({ S3483, S3457 }),
  .out1({ S3486 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3988_ (
  .in1({ S3483, S3457 }),
  .out1({ S3487 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3989_ (
  .in1({ S3484, S3458 }),
  .out1({ S3488 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3990_ (
  .in1({ S3487, S3485 }),
  .out1({ S3490 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3991_ (
  .in1({ S3488, S3486 }),
  .out1({ S3491 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3992_ (
  .in1({ S3491, S3438 }),
  .out1({ S3492 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3993_ (
  .in1({ S3490, S3439 }),
  .out1({ S3493 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3994_ (
  .in1({ S3490, S3439 }),
  .out1({ S3494 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3995_ (
  .in1({ S3491, S3438 }),
  .out1({ S3495 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3996_ (
  .in1({ S3494, S3492 }),
  .out1({ S3496 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3997_ (
  .in1({ S3495, S3493 }),
  .out1({ S3497 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_3998_ (
  .in1({ S3497, S3437 }),
  .out1({ S3498 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_3999_ (
  .in1({ S3496, S3436 }),
  .out1({ S3499 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4000_ (
  .in1({ S3496, S3436 }),
  .out1({ S3501 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4001_ (
  .in1({ S3497, S3437 }),
  .out1({ S3502 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4002_ (
  .in1({ S3501, S3498 }),
  .out1({ S3503 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4003_ (
  .in1({ S3502, S3499 }),
  .out1({ S3504 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4004_ (
  .in1({ S3504, S3398 }),
  .out1({ S3505 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4005_ (
  .in1({ S3503, S3399 }),
  .out1({ S3506 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4006_ (
  .in1({ S3503, S3399 }),
  .out1({ S3507 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4007_ (
  .in1({ S3504, S3398 }),
  .out1({ S3508 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4008_ (
  .in1({ S3507, S3505 }),
  .out1({ S3509 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4009_ (
  .in1({ S3508, S3506 }),
  .out1({ S3510 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4010_ (
  .in1({ S3510, S3397 }),
  .out1({ S3512 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4011_ (
  .in1({ S3509, S3396 }),
  .out1({ S3513 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4012_ (
  .in1({ S3509, S3396 }),
  .out1({ S3514 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4013_ (
  .in1({ S3510, S3397 }),
  .out1({ S3515 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4014_ (
  .in1({ S3514, S3512 }),
  .out1({ S3516 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4015_ (
  .in1({ S3515, S3513 }),
  .out1({ S3517 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4016_ (
  .in1({ S3517, S3348 }),
  .out1({ S3518 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4017_ (
  .in1({ S3516, S3349 }),
  .out1({ S3519 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4018_ (
  .in1({ S3516, S3349 }),
  .out1({ S3520 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4019_ (
  .in1({ S3517, S3348 }),
  .out1({ S3521 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4020_ (
  .in1({ S3520, S3518 }),
  .out1({ S3523 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4021_ (
  .in1({ S3521, S3519 }),
  .out1({ S3524 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4022_ (
  .in1({ S3524, S3196 }),
  .out1({ S3525 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4023_ (
  .in1({ S3523, S3195 }),
  .out1({ S3526 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4024_ (
  .in1({ S3523, S3195 }),
  .out1({ S3527 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4025_ (
  .in1({ S3524, S3196 }),
  .out1({ S3528 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4026_ (
  .in1({ S3527, S3525 }),
  .out1({ S3529 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4027_ (
  .in1({ S3528, S3526 }),
  .out1({ S3530 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4028_ (
  .in1({ S3529, S3347 }),
  .out1({ S3531 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4029_ (
  .in1({ S3530, S3345 }),
  .out1({ S3532 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4030_ (
  .in1({ S3530, S3345 }),
  .out1({ S3534 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4031_ (
  .in1({ S3529, S3347 }),
  .out1({ S3535 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4032_ (
  .in1({ S3534, S3531 }),
  .out1({ S3536 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4033_ (
  .in1({ S3535, S3532 }),
  .out1({ S3537 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4034_ (
  .in1({ S3536, S3332 }),
  .out1({ S3538 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4035_ (
  .in1({ S3537, S3331 }),
  .out1({ S3539 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4036_ (
  .in1({ S3539, S3538 }),
  .out1({ S3540 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4037_ (
  .in1({ S3540, S3344 }),
  .out1({ S3541 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4038_ (
  .in1({ S3541 }),
  .out1({ S3542 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4039_ (
  .in1({ S3540, S3344 }),
  .out1({ S3543 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4040_ (
  .in1({ S3541, S5590 }),
  .out1({ S3545 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4041_ (
  .in1({ S3545, S3543 }),
  .out1({ S3546 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4042_ (
  .in1({ S5611, new_datapath_multdivunit_outmdu1_12 }),
  .out1({ S3547 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4043_ (
  .in1({ S3547 }),
  .out1({ S3548 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4044_ (
  .in1({ S393, S5547 }),
  .out1({ S3549 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4045_ (
  .in1({ S3549, S3548 }),
  .out1({ S3550 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4046_ (
  .in1({ S3550, S3546 }),
  .out1({ S32 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4047_ (
  .in1({ S3542, S3538 }),
  .out1({ S3551 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4048_ (
  .in1({ S3551 }),
  .out1({ S3552 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4049_ (
  .in1({ S3526, S3519 }),
  .out1({ S3553 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4050_ (
  .in1({ S3392, S3385 }),
  .out1({ S3555 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4051_ (
  .in1({ S3393, S3386 }),
  .out1({ S3556 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4052_ (
  .in1({ S3512, S3505 }),
  .out1({ S3557 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4053_ (
  .in1({ S3513, S3506 }),
  .out1({ S3558 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4054_ (
  .in1({ S3376, S3370 }),
  .out1({ S3559 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4055_ (
  .in1({ S3377, S3371 }),
  .out1({ S3560 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4056_ (
  .in1({ new_datapath_addsubunit_in1_0, new_datapath_multdivunit_1697_B_13 }),
  .out1({ S3561 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4057_ (
  .in1({ new_datapath_addsubunit_in1_1, new_datapath_multdivunit_1697_B_12 }),
  .out1({ S3562 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4058_ (
  .in1({ S3562, S3561 }),
  .out1({ S3563 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4059_ (
  .in1({ S3563 }),
  .out1({ S3564 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4060_ (
  .in1({ new_datapath_addsubunit_in1_1, new_datapath_multdivunit_1697_B_13 }),
  .out1({ S3566 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4061_ (
  .in1({ S3566 }),
  .out1({ S3567 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4062_ (
  .in1({ S3566, S3351 }),
  .out1({ S3568 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4063_ (
  .in1({ S3567, S3350 }),
  .out1({ S3569 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4064_ (
  .in1({ S3568, S3564 }),
  .out1({ S3570 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4065_ (
  .in1({ S3569, S3563 }),
  .out1({ S3571 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4066_ (
  .in1({ S3363, S3360 }),
  .out1({ S3572 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4067_ (
  .in1({ S3572 }),
  .out1({ S3573 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4068_ (
  .in1({ new_datapath_addsubunit_in1_2, new_datapath_multdivunit_1697_B_11 }),
  .out1({ S3574 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4069_ (
  .in1({ S3574 }),
  .out1({ S3575 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4070_ (
  .in1({ S5936, S3467 }),
  .out1({ S3577 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4071_ (
  .in1({ new_datapath_addsubunit_in1_4, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S3578 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4072_ (
  .in1({ S3578, S3359 }),
  .out1({ S3579 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4073_ (
  .in1({ new_datapath_addsubunit_in1_4, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S3580 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4074_ (
  .in1({ S3578, S3359 }),
  .out1({ S3581 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4075_ (
  .in1({ S3577, S3358 }),
  .out1({ S3582 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4076_ (
  .in1({ S3582, S3579 }),
  .out1({ S3583 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4077_ (
  .in1({ S3583 }),
  .out1({ S3584 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4078_ (
  .in1({ S3583, S3574 }),
  .out1({ S3585 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4079_ (
  .in1({ S3584, S3575 }),
  .out1({ S3586 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4080_ (
  .in1({ S3583, S3574 }),
  .out1({ S3588 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4081_ (
  .in1({ S3588, S3586 }),
  .out1({ S3589 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4082_ (
  .in1({ S3589 }),
  .out1({ S3590 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4083_ (
  .in1({ S3589, S3572 }),
  .out1({ S3591 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4084_ (
  .in1({ S3590, S3573 }),
  .out1({ S3592 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4085_ (
  .in1({ S3589, S3572 }),
  .out1({ S3593 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4086_ (
  .in1({ S3593 }),
  .out1({ S3594 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4087_ (
  .in1({ S3594, S3591 }),
  .out1({ S3595 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4088_ (
  .in1({ S3593, S3592 }),
  .out1({ S3596 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4089_ (
  .in1({ S3595, S3570 }),
  .out1({ S3597 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4090_ (
  .in1({ S3596, S3571 }),
  .out1({ S3599 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4091_ (
  .in1({ S3596, S3571 }),
  .out1({ S3600 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4092_ (
  .in1({ S3595, S3570 }),
  .out1({ S3601 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4093_ (
  .in1({ S3600, S3597 }),
  .out1({ S3602 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4094_ (
  .in1({ S3601, S3599 }),
  .out1({ S3603 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4095_ (
  .in1({ S3433, S3425 }),
  .out1({ S3604 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4096_ (
  .in1({ S3435, S3426 }),
  .out1({ S3605 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4097_ (
  .in1({ S3604, S3603 }),
  .out1({ S3606 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4098_ (
  .in1({ S3605, S3602 }),
  .out1({ S3607 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4099_ (
  .in1({ S3605, S3602 }),
  .out1({ S3608 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4100_ (
  .in1({ S3604, S3603 }),
  .out1({ S3610 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4101_ (
  .in1({ S3608, S3606 }),
  .out1({ S3611 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4102_ (
  .in1({ S3610, S3607 }),
  .out1({ S3612 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4103_ (
  .in1({ S3611, S3560 }),
  .out1({ S3613 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4104_ (
  .in1({ S3612, S3559 }),
  .out1({ S3614 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4105_ (
  .in1({ S3612, S3559 }),
  .out1({ S3615 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4106_ (
  .in1({ S3611, S3560 }),
  .out1({ S3616 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4107_ (
  .in1({ S3615, S3613 }),
  .out1({ S3617 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4108_ (
  .in1({ S3616, S3614 }),
  .out1({ S3618 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4109_ (
  .in1({ S3498, S3492 }),
  .out1({ S3619 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4110_ (
  .in1({ S3499, S3493 }),
  .out1({ S3621 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4111_ (
  .in1({ S3416, S3411 }),
  .out1({ S3622 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4112_ (
  .in1({ S3417, S3413 }),
  .out1({ S3623 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4113_ (
  .in1({ S5926, S3478 }),
  .out1({ S3624 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4114_ (
  .in1({ new_datapath_addsubunit_in1_5, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S3625 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4115_ (
  .in1({ S202, S5907 }),
  .out1({ S3626 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4116_ (
  .in1({ S203, new_datapath_addsubunit_in1_7 }),
  .out1({ S3627 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4117_ (
  .in1({ S3626, S3409 }),
  .out1({ S3628 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4118_ (
  .in1({ S3627, S3410 }),
  .out1({ S3629 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4119_ (
  .in1({ S229, new_datapath_addsubunit_in1_7 }),
  .out1({ S3630 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4120_ (
  .in1({ S3627, S3410 }),
  .out1({ S3632 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4121_ (
  .in1({ S3626, S3409 }),
  .out1({ S3633 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4122_ (
  .in1({ S3632, S3628 }),
  .out1({ S3634 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4123_ (
  .in1({ S3633, S3629 }),
  .out1({ S3635 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4124_ (
  .in1({ S3635, S3625 }),
  .out1({ S3636 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4125_ (
  .in1({ S3634, S3624 }),
  .out1({ S3637 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4126_ (
  .in1({ S3634, S3624 }),
  .out1({ S3638 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4127_ (
  .in1({ S3635, S3625 }),
  .out1({ S3639 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4128_ (
  .in1({ S3638, S3636 }),
  .out1({ S3640 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4129_ (
  .in1({ S3639, S3637 }),
  .out1({ S3641 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4130_ (
  .in1({ S3452, S3448 }),
  .out1({ S3643 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4131_ (
  .in1({ S3453, S3449 }),
  .out1({ S3644 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4132_ (
  .in1({ S3643, S3641 }),
  .out1({ S3645 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4133_ (
  .in1({ S3644, S3640 }),
  .out1({ S3646 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4134_ (
  .in1({ S3644, S3640 }),
  .out1({ S3647 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4135_ (
  .in1({ S3643, S3641 }),
  .out1({ S3648 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4136_ (
  .in1({ S3647, S3645 }),
  .out1({ S3649 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4137_ (
  .in1({ S3648, S3646 }),
  .out1({ S3650 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4138_ (
  .in1({ S3649, S3623 }),
  .out1({ S3651 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4139_ (
  .in1({ S3650, S3622 }),
  .out1({ S3652 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4140_ (
  .in1({ S3650, S3622 }),
  .out1({ S3654 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4141_ (
  .in1({ S3649, S3623 }),
  .out1({ S3655 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4142_ (
  .in1({ S3654, S3651 }),
  .out1({ S3656 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4143_ (
  .in1({ S3655, S3652 }),
  .out1({ S3657 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4144_ (
  .in1({ S3485, S3479 }),
  .out1({ S3658 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4145_ (
  .in1({ S3486, S3480 }),
  .out1({ S3659 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4146_ (
  .in1({ S209, new_datapath_addsubunit_in1_8 }),
  .out1({ S3660 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4147_ (
  .in1({ S3660 }),
  .out1({ S3661 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4148_ (
  .in1({ S248, S3346 }),
  .out1({ S3662 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4149_ (
  .in1({ S249, new_datapath_addsubunit_in1_10 }),
  .out1({ S3663 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4150_ (
  .in1({ S3663, S3447 }),
  .out1({ S3665 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4151_ (
  .in1({ S241, new_datapath_addsubunit_in1_10 }),
  .out1({ S3666 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4152_ (
  .in1({ S3663, S3447 }),
  .out1({ S3667 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4153_ (
  .in1({ S3662, S3446 }),
  .out1({ S3668 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4154_ (
  .in1({ S3668, S3665 }),
  .out1({ S3669 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4155_ (
  .in1({ S3669 }),
  .out1({ S3670 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4156_ (
  .in1({ S3669, S3660 }),
  .out1({ S3671 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4157_ (
  .in1({ S3670, S3661 }),
  .out1({ S3672 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4158_ (
  .in1({ S3669, S3660 }),
  .out1({ S3673 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4159_ (
  .in1({ S3673 }),
  .out1({ S3674 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4160_ (
  .in1({ S3674, S3671 }),
  .out1({ S3676 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4161_ (
  .in1({ S3673, S3672 }),
  .out1({ S3677 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4162_ (
  .in1({ S3472, S3468 }),
  .out1({ S3678 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4163_ (
  .in1({ S3473, S3469 }),
  .out1({ S3679 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4164_ (
  .in1({ S256, S3357 }),
  .out1({ S3680 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4165_ (
  .in1({ S257, new_datapath_addsubunit_in1_11 }),
  .out1({ S3681 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4166_ (
  .in1({ S3465, S351 }),
  .out1({ S3682 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4167_ (
  .in1({ S3466, S352 }),
  .out1({ S3683 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4168_ (
  .in1({ S265, new_datapath_addsubunit_in1_13 }),
  .out1({ S3684 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4169_ (
  .in1({ S3466, S352 }),
  .out1({ S3685 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4170_ (
  .in1({ S3465, S351 }),
  .out1({ S3687 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4171_ (
  .in1({ S3685, S3682 }),
  .out1({ S3688 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4172_ (
  .in1({ S3687, S3683 }),
  .out1({ S3689 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4173_ (
  .in1({ S3689, S3681 }),
  .out1({ S3690 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4174_ (
  .in1({ S3688, S3680 }),
  .out1({ S3691 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4175_ (
  .in1({ S3688, S3680 }),
  .out1({ S3692 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4176_ (
  .in1({ S3689, S3681 }),
  .out1({ S3693 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4177_ (
  .in1({ S3692, S3690 }),
  .out1({ S3694 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4178_ (
  .in1({ S3693, S3691 }),
  .out1({ S3695 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4179_ (
  .in1({ S3695, S3678 }),
  .out1({ S3696 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4180_ (
  .in1({ S3694, S3679 }),
  .out1({ S3698 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4181_ (
  .in1({ S3694, S3679 }),
  .out1({ S3699 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4182_ (
  .in1({ S3695, S3678 }),
  .out1({ S3700 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4183_ (
  .in1({ S3699, S3696 }),
  .out1({ S3701 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4184_ (
  .in1({ S3700, S3698 }),
  .out1({ S3702 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4185_ (
  .in1({ S3702, S3677 }),
  .out1({ S3703 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4186_ (
  .in1({ S3701, S3676 }),
  .out1({ S3704 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4187_ (
  .in1({ S3701, S3676 }),
  .out1({ S3705 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4188_ (
  .in1({ S3702, S3677 }),
  .out1({ S3706 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4189_ (
  .in1({ S3705, S3703 }),
  .out1({ S3707 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4190_ (
  .in1({ S3706, S3704 }),
  .out1({ S3709 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4191_ (
  .in1({ S3709, S3658 }),
  .out1({ S3710 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4192_ (
  .in1({ S3707, S3659 }),
  .out1({ S3711 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4193_ (
  .in1({ S3707, S3659 }),
  .out1({ S3712 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4194_ (
  .in1({ S3709, S3658 }),
  .out1({ S3713 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4195_ (
  .in1({ S3712, S3710 }),
  .out1({ S3714 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4196_ (
  .in1({ S3713, S3711 }),
  .out1({ S3715 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4197_ (
  .in1({ S3715, S3657 }),
  .out1({ S3716 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4198_ (
  .in1({ S3714, S3656 }),
  .out1({ S3717 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4199_ (
  .in1({ S3714, S3656 }),
  .out1({ S3718 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4200_ (
  .in1({ S3715, S3657 }),
  .out1({ S3720 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4201_ (
  .in1({ S3718, S3716 }),
  .out1({ S3721 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4202_ (
  .in1({ S3720, S3717 }),
  .out1({ S3722 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4203_ (
  .in1({ S3722, S3619 }),
  .out1({ S3723 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4204_ (
  .in1({ S3721, S3621 }),
  .out1({ S3724 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4205_ (
  .in1({ S3721, S3621 }),
  .out1({ S3725 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4206_ (
  .in1({ S3722, S3619 }),
  .out1({ S3726 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4207_ (
  .in1({ S3725, S3723 }),
  .out1({ S3727 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4208_ (
  .in1({ S3726, S3724 }),
  .out1({ S3728 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4209_ (
  .in1({ S3728, S3618 }),
  .out1({ S3729 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4210_ (
  .in1({ S3727, S3617 }),
  .out1({ S3730 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4211_ (
  .in1({ S3727, S3617 }),
  .out1({ S3731 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4212_ (
  .in1({ S3728, S3618 }),
  .out1({ S3732 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4213_ (
  .in1({ S3731, S3729 }),
  .out1({ S3733 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4214_ (
  .in1({ S3732, S3730 }),
  .out1({ S3734 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4215_ (
  .in1({ S3734, S3557 }),
  .out1({ S3735 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4216_ (
  .in1({ S3733, S3558 }),
  .out1({ S3736 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4217_ (
  .in1({ S3733, S3558 }),
  .out1({ S3737 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4218_ (
  .in1({ S3734, S3557 }),
  .out1({ S3738 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4219_ (
  .in1({ S3737, S3735 }),
  .out1({ S3739 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4220_ (
  .in1({ S3738, S3736 }),
  .out1({ S3741 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4221_ (
  .in1({ S3741, S3555 }),
  .out1({ S3742 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4222_ (
  .in1({ S3739, S3556 }),
  .out1({ S3743 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4223_ (
  .in1({ S3743, S3742 }),
  .out1({ S3744 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4224_ (
  .in1({ S3744, S3553 }),
  .out1({ S3745 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4225_ (
  .in1({ S3745 }),
  .out1({ S3746 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4226_ (
  .in1({ S3744, S3553 }),
  .out1({ S3747 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4227_ (
  .in1({ S3747 }),
  .out1({ S3748 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4228_ (
  .in1({ S3748, S3745 }),
  .out1({ S3749 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4229_ (
  .in1({ S3747, S3746 }),
  .out1({ S3750 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4230_ (
  .in1({ S3749, S3534 }),
  .out1({ S3751 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4231_ (
  .in1({ S3750, S3535 }),
  .out1({ S3752 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4232_ (
  .in1({ S3752, S3751 }),
  .out1({ S3753 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4233_ (
  .in1({ S3751, S3552 }),
  .out1({ S3754 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4234_ (
  .in1({ S3753, S3551 }),
  .out1({ S3755 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4235_ (
  .in1({ S3755, S3754 }),
  .out1({ S3756 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4236_ (
  .in1({ S3756, S5579 }),
  .out1({ S3757 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4237_ (
  .in1({ S332, S5547 }),
  .out1({ S3758 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4238_ (
  .in1({ S5611, new_datapath_multdivunit_outmdu1_13 }),
  .out1({ S3759 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4239_ (
  .in1({ S3759 }),
  .out1({ S3760 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4240_ (
  .in1({ S3760, S3758 }),
  .out1({ S3762 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4241_ (
  .in1({ S3762, S3757 }),
  .out1({ S33 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4242_ (
  .in1({ S3742, S3735 }),
  .out1({ S3763 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4243_ (
  .in1({ S3763 }),
  .out1({ S3764 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4244_ (
  .in1({ S3615, S3606 }),
  .out1({ S3765 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4245_ (
  .in1({ S3616, S3607 }),
  .out1({ S3766 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4246_ (
  .in1({ S3765, S3569 }),
  .out1({ S3767 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4247_ (
  .in1({ S3766, S3568 }),
  .out1({ S3768 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4248_ (
  .in1({ S3766, S3568 }),
  .out1({ S3769 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4249_ (
  .in1({ S3765, S3569 }),
  .out1({ S3770 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4250_ (
  .in1({ S3769, S3767 }),
  .out1({ S3772 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4251_ (
  .in1({ S3770, S3768 }),
  .out1({ S3773 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4252_ (
  .in1({ S3729, S3723 }),
  .out1({ S3774 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4253_ (
  .in1({ S3730, S3724 }),
  .out1({ S3775 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4254_ (
  .in1({ S3600, S3591 }),
  .out1({ S3776 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4255_ (
  .in1({ S3601, S3592 }),
  .out1({ S3777 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4256_ (
  .in1({ new_datapath_addsubunit_in1_0, new_datapath_multdivunit_1697_B_14 }),
  .out1({ S3778 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4257_ (
  .in1({ new_datapath_addsubunit_in1_2, new_datapath_multdivunit_1697_B_12 }),
  .out1({ S3779 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4258_ (
  .in1({ S3779, S3566 }),
  .out1({ S3780 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4259_ (
  .in1({ S5957, S3423 }),
  .out1({ S3781 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4260_ (
  .in1({ new_datapath_addsubunit_in1_2, new_datapath_multdivunit_1697_B_13 }),
  .out1({ S3783 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4261_ (
  .in1({ S3783, S3562 }),
  .out1({ S3784 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4262_ (
  .in1({ S3784 }),
  .out1({ S3785 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4263_ (
  .in1({ S3785, S3780 }),
  .out1({ S3786 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4264_ (
  .in1({ S3786, S3778 }),
  .out1({ S3787 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4265_ (
  .in1({ S3787 }),
  .out1({ S3788 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4266_ (
  .in1({ S3786, S3778 }),
  .out1({ S3789 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4267_ (
  .in1({ S3789 }),
  .out1({ S3790 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4268_ (
  .in1({ S3790, S3787 }),
  .out1({ S3791 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4269_ (
  .in1({ S3789, S3788 }),
  .out1({ S3792 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4270_ (
  .in1({ S3585, S3581 }),
  .out1({ S3794 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4271_ (
  .in1({ S3586, S3582 }),
  .out1({ S3795 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4272_ (
  .in1({ new_datapath_addsubunit_in1_3, new_datapath_multdivunit_1697_B_11 }),
  .out1({ S3796 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4273_ (
  .in1({ S3796 }),
  .out1({ S3797 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4274_ (
  .in1({ new_datapath_addsubunit_in1_5, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S3798 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4275_ (
  .in1({ S3798, S3580 }),
  .out1({ S3799 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4276_ (
  .in1({ S5926, S3456 }),
  .out1({ S3800 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4277_ (
  .in1({ new_datapath_addsubunit_in1_5, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S3801 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4278_ (
  .in1({ S3801, S3578 }),
  .out1({ S3802 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4279_ (
  .in1({ S3800, S3577 }),
  .out1({ S3803 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4280_ (
  .in1({ S3803, S3799 }),
  .out1({ S3805 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4281_ (
  .in1({ S3805 }),
  .out1({ S3806 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4282_ (
  .in1({ S3805, S3796 }),
  .out1({ S3807 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4283_ (
  .in1({ S3806, S3797 }),
  .out1({ S3808 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4284_ (
  .in1({ S3805, S3796 }),
  .out1({ S3809 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4285_ (
  .in1({ S3809 }),
  .out1({ S3810 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4286_ (
  .in1({ S3810, S3807 }),
  .out1({ S3811 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4287_ (
  .in1({ S3809, S3808 }),
  .out1({ S3812 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4288_ (
  .in1({ S3812, S3794 }),
  .out1({ S3813 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4289_ (
  .in1({ S3811, S3795 }),
  .out1({ S3814 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4290_ (
  .in1({ S3811, S3795 }),
  .out1({ S3816 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4291_ (
  .in1({ S3812, S3794 }),
  .out1({ S3817 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4292_ (
  .in1({ S3816, S3813 }),
  .out1({ S3818 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4293_ (
  .in1({ S3817, S3814 }),
  .out1({ S3819 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4294_ (
  .in1({ S3818, S3791 }),
  .out1({ S3820 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4295_ (
  .in1({ S3819, S3792 }),
  .out1({ S3821 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4296_ (
  .in1({ S3819, S3792 }),
  .out1({ S3822 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4297_ (
  .in1({ S3818, S3791 }),
  .out1({ S3823 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4298_ (
  .in1({ S3822, S3820 }),
  .out1({ S3824 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4299_ (
  .in1({ S3823, S3821 }),
  .out1({ S3825 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4300_ (
  .in1({ S3654, S3645 }),
  .out1({ S3827 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4301_ (
  .in1({ S3655, S3646 }),
  .out1({ S3828 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4302_ (
  .in1({ S3827, S3825 }),
  .out1({ S3829 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4303_ (
  .in1({ S3828, S3824 }),
  .out1({ S3830 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4304_ (
  .in1({ S3828, S3824 }),
  .out1({ S3831 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4305_ (
  .in1({ S3827, S3825 }),
  .out1({ S3832 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4306_ (
  .in1({ S3831, S3829 }),
  .out1({ S3833 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4307_ (
  .in1({ S3832, S3830 }),
  .out1({ S3834 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4308_ (
  .in1({ S3833, S3777 }),
  .out1({ S3835 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4309_ (
  .in1({ S3834, S3776 }),
  .out1({ S3836 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4310_ (
  .in1({ S3834, S3776 }),
  .out1({ S3838 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4311_ (
  .in1({ S3833, S3777 }),
  .out1({ S3839 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4312_ (
  .in1({ S3838, S3835 }),
  .out1({ S3840 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4313_ (
  .in1({ S3839, S3836 }),
  .out1({ S3841 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4314_ (
  .in1({ S3716, S3710 }),
  .out1({ S3842 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4315_ (
  .in1({ S3717, S3711 }),
  .out1({ S3843 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4316_ (
  .in1({ S3636, S3632 }),
  .out1({ S3844 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4317_ (
  .in1({ S3637, S3633 }),
  .out1({ S3845 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4318_ (
  .in1({ new_datapath_addsubunit_in1_6, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S3846 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4319_ (
  .in1({ S3846 }),
  .out1({ S3847 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4320_ (
  .in1({ S203, new_datapath_addsubunit_in1_8 }),
  .out1({ S3849 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4321_ (
  .in1({ S3849, S3630 }),
  .out1({ S3850 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4322_ (
  .in1({ S228, S3325 }),
  .out1({ S3851 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4323_ (
  .in1({ S229, new_datapath_addsubunit_in1_8 }),
  .out1({ S3852 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4324_ (
  .in1({ S3852, S3627 }),
  .out1({ S3853 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4325_ (
  .in1({ S3851, S3626 }),
  .out1({ S3854 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4326_ (
  .in1({ S3854, S3850 }),
  .out1({ S3855 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4327_ (
  .in1({ S3855 }),
  .out1({ S3856 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4328_ (
  .in1({ S3855, S3846 }),
  .out1({ S3857 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4329_ (
  .in1({ S3856, S3847 }),
  .out1({ S3858 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4330_ (
  .in1({ S3855, S3846 }),
  .out1({ S3860 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4331_ (
  .in1({ S3860 }),
  .out1({ S3861 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4332_ (
  .in1({ S3861, S3857 }),
  .out1({ S3862 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4333_ (
  .in1({ S3860, S3858 }),
  .out1({ S3863 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4334_ (
  .in1({ S3671, S3667 }),
  .out1({ S3864 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4335_ (
  .in1({ S3672, S3668 }),
  .out1({ S3865 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4336_ (
  .in1({ S3864, S3863 }),
  .out1({ S3866 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4337_ (
  .in1({ S3865, S3862 }),
  .out1({ S3867 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4338_ (
  .in1({ S3865, S3862 }),
  .out1({ S3868 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4339_ (
  .in1({ S3864, S3863 }),
  .out1({ S3869 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4340_ (
  .in1({ S3868, S3866 }),
  .out1({ S3871 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4341_ (
  .in1({ S3869, S3867 }),
  .out1({ S3872 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4342_ (
  .in1({ S3871, S3845 }),
  .out1({ S3873 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4343_ (
  .in1({ S3872, S3844 }),
  .out1({ S3874 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4344_ (
  .in1({ S3872, S3844 }),
  .out1({ S3875 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4345_ (
  .in1({ S3871, S3845 }),
  .out1({ S3876 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4346_ (
  .in1({ S3875, S3873 }),
  .out1({ S3877 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4347_ (
  .in1({ S3876, S3874 }),
  .out1({ S3878 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4348_ (
  .in1({ S3703, S3696 }),
  .out1({ S3879 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4349_ (
  .in1({ S3704, S3698 }),
  .out1({ S3880 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4350_ (
  .in1({ S209, new_datapath_addsubunit_in1_9 }),
  .out1({ S3882 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4351_ (
  .in1({ S3882 }),
  .out1({ S3883 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4352_ (
  .in1({ S249, new_datapath_addsubunit_in1_11 }),
  .out1({ S3884 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4353_ (
  .in1({ S3884, S3666 }),
  .out1({ S3885 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4354_ (
  .in1({ S240, S3357 }),
  .out1({ S3886 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4355_ (
  .in1({ S241, new_datapath_addsubunit_in1_11 }),
  .out1({ S3887 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4356_ (
  .in1({ S3887, S3663 }),
  .out1({ S3888 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4357_ (
  .in1({ S3886, S3662 }),
  .out1({ S3889 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4358_ (
  .in1({ S3889, S3885 }),
  .out1({ S3890 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4359_ (
  .in1({ S3890 }),
  .out1({ S3891 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4360_ (
  .in1({ S3890, S3882 }),
  .out1({ S3893 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4361_ (
  .in1({ S3891, S3883 }),
  .out1({ S3894 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4362_ (
  .in1({ S3890, S3882 }),
  .out1({ S3895 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4363_ (
  .in1({ S3895 }),
  .out1({ S3896 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4364_ (
  .in1({ S3896, S3893 }),
  .out1({ S3897 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4365_ (
  .in1({ S3895, S3894 }),
  .out1({ S3898 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4366_ (
  .in1({ S3690, S3685 }),
  .out1({ S3899 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4367_ (
  .in1({ S3691, S3687 }),
  .out1({ S3900 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4368_ (
  .in1({ S257, new_datapath_addsubunit_in1_12 }),
  .out1({ S3901 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4369_ (
  .in1({ S3901 }),
  .out1({ S3902 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4370_ (
  .in1({ S271, new_datapath_addsubunit_in1_14 }),
  .out1({ S3904 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4371_ (
  .in1({ S3904, S3684 }),
  .out1({ S3905 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4372_ (
  .in1({ S264, S3390 }),
  .out1({ S3906 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4373_ (
  .in1({ S265, new_datapath_addsubunit_in1_14 }),
  .out1({ S3907 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4374_ (
  .in1({ S3907, S352 }),
  .out1({ S3908 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4375_ (
  .in1({ S3906, S351 }),
  .out1({ S3909 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4376_ (
  .in1({ S3909, S3905 }),
  .out1({ S3910 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4377_ (
  .in1({ S3910 }),
  .out1({ S3911 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4378_ (
  .in1({ S3910, S3901 }),
  .out1({ S3912 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4379_ (
  .in1({ S3911, S3902 }),
  .out1({ S3913 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4380_ (
  .in1({ S3910, S3901 }),
  .out1({ S3915 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4381_ (
  .in1({ S3915 }),
  .out1({ S3916 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4382_ (
  .in1({ S3916, S3912 }),
  .out1({ S3917 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4383_ (
  .in1({ S3915, S3913 }),
  .out1({ S3918 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4384_ (
  .in1({ S3918, S3899 }),
  .out1({ S3919 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4385_ (
  .in1({ S3917, S3900 }),
  .out1({ S3920 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4386_ (
  .in1({ S3917, S3900 }),
  .out1({ S3921 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4387_ (
  .in1({ S3918, S3899 }),
  .out1({ S3922 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4388_ (
  .in1({ S3921, S3919 }),
  .out1({ S3923 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4389_ (
  .in1({ S3922, S3920 }),
  .out1({ S3924 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4390_ (
  .in1({ S3924, S3898 }),
  .out1({ S3926 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4391_ (
  .in1({ S3923, S3897 }),
  .out1({ S3927 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4392_ (
  .in1({ S3923, S3897 }),
  .out1({ S3928 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4393_ (
  .in1({ S3924, S3898 }),
  .out1({ S3929 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4394_ (
  .in1({ S3928, S3926 }),
  .out1({ S3930 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4395_ (
  .in1({ S3929, S3927 }),
  .out1({ S3931 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4396_ (
  .in1({ S3931, S3879 }),
  .out1({ S3932 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4397_ (
  .in1({ S3930, S3880 }),
  .out1({ S3933 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4398_ (
  .in1({ S3930, S3880 }),
  .out1({ S3934 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4399_ (
  .in1({ S3931, S3879 }),
  .out1({ S3935 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4400_ (
  .in1({ S3934, S3932 }),
  .out1({ S3937 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4401_ (
  .in1({ S3935, S3933 }),
  .out1({ S3938 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4402_ (
  .in1({ S3938, S3878 }),
  .out1({ S3939 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4403_ (
  .in1({ S3937, S3877 }),
  .out1({ S3940 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4404_ (
  .in1({ S3937, S3877 }),
  .out1({ S3941 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4405_ (
  .in1({ S3938, S3878 }),
  .out1({ S3942 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4406_ (
  .in1({ S3941, S3939 }),
  .out1({ S3943 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4407_ (
  .in1({ S3942, S3940 }),
  .out1({ S3944 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4408_ (
  .in1({ S3944, S3842 }),
  .out1({ S3945 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4409_ (
  .in1({ S3943, S3843 }),
  .out1({ S3946 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4410_ (
  .in1({ S3943, S3843 }),
  .out1({ S3948 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4411_ (
  .in1({ S3944, S3842 }),
  .out1({ S3949 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4412_ (
  .in1({ S3948, S3945 }),
  .out1({ S3950 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4413_ (
  .in1({ S3949, S3946 }),
  .out1({ S3951 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4414_ (
  .in1({ S3951, S3841 }),
  .out1({ S3952 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4415_ (
  .in1({ S3950, S3840 }),
  .out1({ S3953 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4416_ (
  .in1({ S3950, S3840 }),
  .out1({ S3954 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4417_ (
  .in1({ S3951, S3841 }),
  .out1({ S3955 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4418_ (
  .in1({ S3954, S3952 }),
  .out1({ S3956 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4419_ (
  .in1({ S3955, S3953 }),
  .out1({ S3957 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4420_ (
  .in1({ S3957, S3774 }),
  .out1({ S3959 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4421_ (
  .in1({ S3956, S3775 }),
  .out1({ S3960 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4422_ (
  .in1({ S3956, S3775 }),
  .out1({ S3961 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4423_ (
  .in1({ S3957, S3774 }),
  .out1({ S3962 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4424_ (
  .in1({ S3961, S3959 }),
  .out1({ S3963 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4425_ (
  .in1({ S3962, S3960 }),
  .out1({ S3964 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4426_ (
  .in1({ S3964, S3773 }),
  .out1({ S3965 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4427_ (
  .in1({ S3963, S3772 }),
  .out1({ S3966 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4428_ (
  .in1({ S3964, S3773 }),
  .out1({ S3967 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4429_ (
  .in1({ S3967, S3966 }),
  .out1({ S3968 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4430_ (
  .in1({ S3968 }),
  .out1({ S3970 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4431_ (
  .in1({ S3968, S3763 }),
  .out1({ S3971 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4432_ (
  .in1({ S3970, S3764 }),
  .out1({ S3972 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4433_ (
  .in1({ S3972, S3971 }),
  .out1({ S3973 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4434_ (
  .in1({ S3973, S3747 }),
  .out1({ S3974 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4435_ (
  .in1({ S3974 }),
  .out1({ S3975 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4436_ (
  .in1({ S3973, S3747 }),
  .out1({ S3976 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4437_ (
  .in1({ S3976, S3975 }),
  .out1({ S3977 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4438_ (
  .in1({ S3754, S3752 }),
  .out1({ S3978 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4439_ (
  .in1({ S3978, S3977 }),
  .out1({ S3979 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4440_ (
  .in1({ S3978, S3977 }),
  .out1({ S3981 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4441_ (
  .in1({ S3979, S5590 }),
  .out1({ S3982 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4442_ (
  .in1({ S3982, S3981 }),
  .out1({ S3983 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4443_ (
  .in1({ S5611, new_datapath_multdivunit_outmdu1_14 }),
  .out1({ S3984 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4444_ (
  .in1({ S3984 }),
  .out1({ S3985 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4445_ (
  .in1({ S291, S5547 }),
  .out1({ S3986 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4446_ (
  .in1({ S3986, S3985 }),
  .out1({ S3987 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4447_ (
  .in1({ S3987, S3983 }),
  .out1({ S34 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4448_ (
  .in1({ S3979, S3974 }),
  .out1({ S3988 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4449_ (
  .in1({ S3965, S3959 }),
  .out1({ S3989 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4450_ (
  .in1({ S3966, S3960 }),
  .out1({ S3991 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4451_ (
  .in1({ S3822, S3813 }),
  .out1({ S3992 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4452_ (
  .in1({ S3823, S3814 }),
  .out1({ S3993 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4453_ (
  .in1({ S3939, S3932 }),
  .out1({ S3994 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4454_ (
  .in1({ S3940, S3933 }),
  .out1({ S3995 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4455_ (
  .in1({ S3995, S3992 }),
  .out1({ S3996 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4456_ (
  .in1({ S3994, S3993 }),
  .out1({ S3997 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4457_ (
  .in1({ S3994, S3993 }),
  .out1({ S3998 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4458_ (
  .in1({ S3995, S3992 }),
  .out1({ S3999 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4459_ (
  .in1({ S3998, S3996 }),
  .out1({ S4000 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4460_ (
  .in1({ S3999, S3997 }),
  .out1({ S4002 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4461_ (
  .in1({ S3952, S3945 }),
  .out1({ S4003 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4462_ (
  .in1({ S3953, S3946 }),
  .out1({ S4004 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4463_ (
  .in1({ S3875, S3866 }),
  .out1({ S4005 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4464_ (
  .in1({ S3876, S3867 }),
  .out1({ S4006 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4465_ (
  .in1({ S3807, S3802 }),
  .out1({ S4007 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4466_ (
  .in1({ S3808, S3803 }),
  .out1({ S4008 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4467_ (
  .in1({ S5936, S3445 }),
  .out1({ S4009 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4468_ (
  .in1({ new_datapath_addsubunit_in1_4, new_datapath_multdivunit_1697_B_11 }),
  .out1({ S4010 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4469_ (
  .in1({ S5916, S3467 }),
  .out1({ S4011 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4470_ (
  .in1({ new_datapath_addsubunit_in1_6, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S4013 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4471_ (
  .in1({ S4013, S3800 }),
  .out1({ S4014 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4472_ (
  .in1({ S4011, S3801 }),
  .out1({ S4015 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4473_ (
  .in1({ S4011, S3801 }),
  .out1({ S4016 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4474_ (
  .in1({ S4013, S3800 }),
  .out1({ S4017 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4475_ (
  .in1({ S4016, S4014 }),
  .out1({ S4018 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4476_ (
  .in1({ S4017, S4015 }),
  .out1({ S4019 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4477_ (
  .in1({ S4019, S4010 }),
  .out1({ S4020 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4478_ (
  .in1({ S4018, S4009 }),
  .out1({ S4021 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4479_ (
  .in1({ S4018, S4009 }),
  .out1({ S4022 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4480_ (
  .in1({ S4019, S4010 }),
  .out1({ S4024 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4481_ (
  .in1({ S4022, S4020 }),
  .out1({ S4025 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4482_ (
  .in1({ S4024, S4021 }),
  .out1({ S4026 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4483_ (
  .in1({ S4026, S4007 }),
  .out1({ S4027 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4484_ (
  .in1({ S4025, S4008 }),
  .out1({ S4028 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4485_ (
  .in1({ S4025, S4008 }),
  .out1({ S4029 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4486_ (
  .in1({ S4026, S4007 }),
  .out1({ S4030 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4487_ (
  .in1({ S4029, S4027 }),
  .out1({ S4031 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4488_ (
  .in1({ S4030, S4028 }),
  .out1({ S4032 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4489_ (
  .in1({ S4032, S4006 }),
  .out1({ S4033 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4490_ (
  .in1({ S4031, S4005 }),
  .out1({ S4035 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4491_ (
  .in1({ S4031, S4005 }),
  .out1({ S4036 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4492_ (
  .in1({ S4032, S4006 }),
  .out1({ S4037 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4493_ (
  .in1({ S4036, S4033 }),
  .out1({ S4038 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4494_ (
  .in1({ S4037, S4035 }),
  .out1({ S4039 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4495_ (
  .in1({ S248, S3368 }),
  .out1({ S4040 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4496_ (
  .in1({ S249, new_datapath_addsubunit_in1_12 }),
  .out1({ S4041 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4497_ (
  .in1({ S270, S3401 }),
  .out1({ S4042 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4498_ (
  .in1({ S271, new_datapath_addsubunit_in1_15 }),
  .out1({ S4043 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4499_ (
  .in1({ S4043, S3906 }),
  .out1({ S4044 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4500_ (
  .in1({ S4042, S3907 }),
  .out1({ S4046 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4501_ (
  .in1({ S4042, S3907 }),
  .out1({ S4047 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4502_ (
  .in1({ S4043, S3906 }),
  .out1({ S4048 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4503_ (
  .in1({ S4047, S4044 }),
  .out1({ S4049 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4504_ (
  .in1({ S4048, S4046 }),
  .out1({ S4050 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4505_ (
  .in1({ S208, S3346 }),
  .out1({ S4051 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4506_ (
  .in1({ S209, new_datapath_addsubunit_in1_10 }),
  .out1({ S4052 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4507_ (
  .in1({ S256, S3379 }),
  .out1({ S4053 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4508_ (
  .in1({ S257, new_datapath_addsubunit_in1_13 }),
  .out1({ S4054 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4509_ (
  .in1({ S3912, S3908 }),
  .out1({ S4055 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4510_ (
  .in1({ S3913, S3909 }),
  .out1({ S4057 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4511_ (
  .in1({ S4041, S3886 }),
  .out1({ S4058 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4512_ (
  .in1({ S4040, S3887 }),
  .out1({ S4059 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4513_ (
  .in1({ S4040, S3887 }),
  .out1({ S4060 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4514_ (
  .in1({ S4041, S3886 }),
  .out1({ S4061 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4515_ (
  .in1({ S4060, S4058 }),
  .out1({ S4062 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4516_ (
  .in1({ S4061, S4059 }),
  .out1({ S4063 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4517_ (
  .in1({ S4063, S4052 }),
  .out1({ S4064 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4518_ (
  .in1({ S4062, S4051 }),
  .out1({ S4065 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4519_ (
  .in1({ S4062, S4051 }),
  .out1({ S4066 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4520_ (
  .in1({ S4063, S4052 }),
  .out1({ S4068 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4521_ (
  .in1({ S4066, S4064 }),
  .out1({ S4069 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4522_ (
  .in1({ S4068, S4065 }),
  .out1({ S4070 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4523_ (
  .in1({ S4054, S4050 }),
  .out1({ S4071 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4524_ (
  .in1({ S4053, S4049 }),
  .out1({ S4072 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4525_ (
  .in1({ S4053, S4049 }),
  .out1({ S4073 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4526_ (
  .in1({ S4054, S4050 }),
  .out1({ S4074 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4527_ (
  .in1({ S4073, S4071 }),
  .out1({ S4075 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4528_ (
  .in1({ S4074, S4072 }),
  .out1({ S4076 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4529_ (
  .in1({ S4075, S4055 }),
  .out1({ S4077 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4530_ (
  .in1({ S4076, S4057 }),
  .out1({ S4079 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4531_ (
  .in1({ S4076, S4057 }),
  .out1({ S4080 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4532_ (
  .in1({ S4075, S4055 }),
  .out1({ S4081 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4533_ (
  .in1({ S4080, S4077 }),
  .out1({ S4082 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4534_ (
  .in1({ S4081, S4079 }),
  .out1({ S4083 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4535_ (
  .in1({ S4083, S4069 }),
  .out1({ S4084 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4536_ (
  .in1({ S4082, S4070 }),
  .out1({ S4085 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4537_ (
  .in1({ S4082, S4070 }),
  .out1({ S4086 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4538_ (
  .in1({ S4083, S4069 }),
  .out1({ S4087 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4539_ (
  .in1({ S4086, S4084 }),
  .out1({ S4088 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4540_ (
  .in1({ S4087, S4085 }),
  .out1({ S4090 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4541_ (
  .in1({ S5907, S3478 }),
  .out1({ S4091 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4542_ (
  .in1({ new_datapath_addsubunit_in1_7, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S4092 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4543_ (
  .in1({ S3893, S3888 }),
  .out1({ S4093 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4544_ (
  .in1({ S3894, S3889 }),
  .out1({ S4094 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4545_ (
  .in1({ S202, S3336 }),
  .out1({ S4095 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4546_ (
  .in1({ S203, new_datapath_addsubunit_in1_9 }),
  .out1({ S4096 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4547_ (
  .in1({ S4096, S3851 }),
  .out1({ S4097 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4548_ (
  .in1({ S4095, S3852 }),
  .out1({ S4098 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4549_ (
  .in1({ S4095, S3852 }),
  .out1({ S4099 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4550_ (
  .in1({ S4096, S3851 }),
  .out1({ S4101 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4551_ (
  .in1({ S4099, S4097 }),
  .out1({ S4102 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4552_ (
  .in1({ S4101, S4098 }),
  .out1({ S4103 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4553_ (
  .in1({ S4103, S4094 }),
  .out1({ S4104 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4554_ (
  .in1({ S4102, S4093 }),
  .out1({ S4105 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4555_ (
  .in1({ S4102, S4093 }),
  .out1({ S4106 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4556_ (
  .in1({ S4103, S4094 }),
  .out1({ S4107 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4557_ (
  .in1({ S4106, S4104 }),
  .out1({ S4108 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4558_ (
  .in1({ S4107, S4105 }),
  .out1({ S4109 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4559_ (
  .in1({ S4109, S4091 }),
  .out1({ S4110 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4560_ (
  .in1({ S4108, S4092 }),
  .out1({ S4112 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4561_ (
  .in1({ S4108, S4092 }),
  .out1({ S4113 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4562_ (
  .in1({ S4109, S4091 }),
  .out1({ S4114 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4563_ (
  .in1({ S4113, S4110 }),
  .out1({ S4115 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4564_ (
  .in1({ S4114, S4112 }),
  .out1({ S4116 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4565_ (
  .in1({ S4116, S4090 }),
  .out1({ S4117 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4566_ (
  .in1({ S4115, S4088 }),
  .out1({ S4118 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4567_ (
  .in1({ S4115, S4088 }),
  .out1({ S4119 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4568_ (
  .in1({ S4116, S4090 }),
  .out1({ S4120 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4569_ (
  .in1({ S4119, S4117 }),
  .out1({ S4121 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4570_ (
  .in1({ S4120, S4118 }),
  .out1({ S4123 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4571_ (
  .in1({ new_datapath_addsubunit_in1_0, new_datapath_multdivunit_1697_B_15 }),
  .out1({ S4124 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4572_ (
  .in1({ S5966, S3412 }),
  .out1({ S4125 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4573_ (
  .in1({ new_datapath_addsubunit_in1_1, new_datapath_multdivunit_1697_B_14 }),
  .out1({ S4126 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4574_ (
  .in1({ S5947, S3434 }),
  .out1({ S4127 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4575_ (
  .in1({ new_datapath_addsubunit_in1_3, new_datapath_multdivunit_1697_B_12 }),
  .out1({ S4128 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4576_ (
  .in1({ S4128, S3781 }),
  .out1({ S4129 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4577_ (
  .in1({ S4127, S3783 }),
  .out1({ S4130 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4578_ (
  .in1({ S4127, S3783 }),
  .out1({ S4131 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4579_ (
  .in1({ S4128, S3781 }),
  .out1({ S4132 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4580_ (
  .in1({ S4131, S4129 }),
  .out1({ S4134 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4581_ (
  .in1({ S4132, S4130 }),
  .out1({ S4135 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4582_ (
  .in1({ S4135, S4126 }),
  .out1({ S4136 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4583_ (
  .in1({ S4134, S4125 }),
  .out1({ S4137 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4584_ (
  .in1({ S4134, S4125 }),
  .out1({ S4138 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4585_ (
  .in1({ S4135, S4126 }),
  .out1({ S4139 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4586_ (
  .in1({ S4138, S4136 }),
  .out1({ S4140 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4587_ (
  .in1({ S4139, S4137 }),
  .out1({ S4141 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4588_ (
  .in1({ S3787, S3784 }),
  .out1({ S4142 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4589_ (
  .in1({ S3857, S3853 }),
  .out1({ S4143 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4590_ (
  .in1({ S3858, S3854 }),
  .out1({ S4145 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4591_ (
  .in1({ S3926, S3919 }),
  .out1({ S4146 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4592_ (
  .in1({ S3927, S3920 }),
  .out1({ S4147 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4593_ (
  .in1({ S4147, S4143 }),
  .out1({ S4148 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4594_ (
  .in1({ S4146, S4145 }),
  .out1({ S4149 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4595_ (
  .in1({ S4146, S4145 }),
  .out1({ S4150 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4596_ (
  .in1({ S4147, S4143 }),
  .out1({ S4151 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4597_ (
  .in1({ S4150, S4148 }),
  .out1({ S4152 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4598_ (
  .in1({ S4151, S4149 }),
  .out1({ S4153 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4599_ (
  .in1({ S4153, S4123 }),
  .out1({ S4154 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4600_ (
  .in1({ S4152, S4121 }),
  .out1({ S4156 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4601_ (
  .in1({ S4152, S4121 }),
  .out1({ S4157 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4602_ (
  .in1({ S4153, S4123 }),
  .out1({ S4158 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4603_ (
  .in1({ S4157, S4154 }),
  .out1({ S4159 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4604_ (
  .in1({ S4158, S4156 }),
  .out1({ S4160 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4605_ (
  .in1({ S4142, S4124 }),
  .out1({ S4161 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4606_ (
  .in1({ S4161 }),
  .out1({ S4162 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4607_ (
  .in1({ S4142, S4124 }),
  .out1({ S4163 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4608_ (
  .in1({ S4163 }),
  .out1({ S4164 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4609_ (
  .in1({ S4163, S4162 }),
  .out1({ S4165 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4610_ (
  .in1({ S4164, S4161 }),
  .out1({ S4167 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4611_ (
  .in1({ S4167, S4140 }),
  .out1({ S4168 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4612_ (
  .in1({ S4165, S4141 }),
  .out1({ S4169 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4613_ (
  .in1({ S4165, S4141 }),
  .out1({ S4170 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4614_ (
  .in1({ S4167, S4140 }),
  .out1({ S4171 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4615_ (
  .in1({ S4170, S4168 }),
  .out1({ S4172 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4616_ (
  .in1({ S4171, S4169 }),
  .out1({ S4173 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4617_ (
  .in1({ S4172, S4160 }),
  .out1({ S4174 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4618_ (
  .in1({ S4173, S4159 }),
  .out1({ S4175 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4619_ (
  .in1({ S4173, S4159 }),
  .out1({ S4176 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4620_ (
  .in1({ S4172, S4160 }),
  .out1({ S4178 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4621_ (
  .in1({ S4176, S4174 }),
  .out1({ S4179 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4622_ (
  .in1({ S4178, S4175 }),
  .out1({ S4180 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4623_ (
  .in1({ S4180, S4039 }),
  .out1({ S4181 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4624_ (
  .in1({ S4179, S4038 }),
  .out1({ S4182 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4625_ (
  .in1({ S4179, S4038 }),
  .out1({ S4183 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4626_ (
  .in1({ S4180, S4039 }),
  .out1({ S4184 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4627_ (
  .in1({ S4183, S4181 }),
  .out1({ S4185 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4628_ (
  .in1({ S4184, S4182 }),
  .out1({ S4186 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4629_ (
  .in1({ S3838, S3829 }),
  .out1({ S4187 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4630_ (
  .in1({ S3839, S3830 }),
  .out1({ S4189 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4631_ (
  .in1({ S4187, S4186 }),
  .out1({ S4190 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4632_ (
  .in1({ S4189, S4185 }),
  .out1({ S4191 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4633_ (
  .in1({ S4189, S4185 }),
  .out1({ S4192 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4634_ (
  .in1({ S4187, S4186 }),
  .out1({ S4193 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4635_ (
  .in1({ S4192, S4190 }),
  .out1({ S4194 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4636_ (
  .in1({ S4193, S4191 }),
  .out1({ S4195 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4637_ (
  .in1({ S4194, S4004 }),
  .out1({ S4196 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4638_ (
  .in1({ S4195, S4003 }),
  .out1({ S4197 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4639_ (
  .in1({ S4195, S4003 }),
  .out1({ S4198 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4640_ (
  .in1({ S4194, S4004 }),
  .out1({ S4200 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4641_ (
  .in1({ S4198, S4196 }),
  .out1({ S4201 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4642_ (
  .in1({ S4200, S4197 }),
  .out1({ S4202 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4643_ (
  .in1({ S4201, S4000 }),
  .out1({ S4203 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4644_ (
  .in1({ S4202, S4002 }),
  .out1({ S4204 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4645_ (
  .in1({ S4202, S4002 }),
  .out1({ S4205 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4646_ (
  .in1({ S4201, S4000 }),
  .out1({ S4206 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4647_ (
  .in1({ S4205, S4203 }),
  .out1({ S4207 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4648_ (
  .in1({ S4206, S4204 }),
  .out1({ S4208 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4649_ (
  .in1({ S4208, S3989 }),
  .out1({ S4209 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4650_ (
  .in1({ S4207, S3991 }),
  .out1({ S4211 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4651_ (
  .in1({ S4207, S3991 }),
  .out1({ S4212 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4652_ (
  .in1({ S4208, S3989 }),
  .out1({ S4213 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4653_ (
  .in1({ S4212, S4209 }),
  .out1({ S4214 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4654_ (
  .in1({ S4213, S4211 }),
  .out1({ S4215 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4655_ (
  .in1({ S3972, S3768 }),
  .out1({ S4216 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4656_ (
  .in1({ S4216 }),
  .out1({ S4217 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4657_ (
  .in1({ S3972, S3768 }),
  .out1({ S4218 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4658_ (
  .in1({ S4218 }),
  .out1({ S4219 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4659_ (
  .in1({ S4218, S4217 }),
  .out1({ S4220 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4660_ (
  .in1({ S4219, S4216 }),
  .out1({ S4222 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4661_ (
  .in1({ S4222, S4214 }),
  .out1({ S4223 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4662_ (
  .in1({ S4220, S4215 }),
  .out1({ S4224 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4663_ (
  .in1({ S4224, S4223 }),
  .out1({ S4225 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4664_ (
  .in1({ S4225, S3988 }),
  .out1({ S4226 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4665_ (
  .in1({ S4225, S3988 }),
  .out1({ S4227 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4666_ (
  .in1({ S4227, S5579 }),
  .out1({ S4228 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4667_ (
  .in1({ S4228, S4226 }),
  .out1({ S4229 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4668_ (
  .in1({ S5611, new_datapath_multdivunit_outmdu1_15 }),
  .out1({ S4230 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4669_ (
  .in1({ S270, new_datapath_addsubunit_in1_15 }),
  .out1({ S4231 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4670_ (
  .in1({ S4231, S5547 }),
  .out1({ S4233 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4671_ (
  .in1({ S4233, S272 }),
  .out1({ S4234 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4672_ (
  .in1({ S4234, S4230 }),
  .out1({ S4235 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4673_ (
  .in1({ S4235, S4229 }),
  .out1({ S4236 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4674_ (
  .in1({ S4236 }),
  .out1({ S35 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4675_ (
  .in1({ S6086, S2800 }),
  .out1({ S36 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4676_ (
  .in1({ S6086, S2811 }),
  .out1({ S37 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4677_ (
  .in1({ S6086, S2822 }),
  .out1({ S38 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4678_ (
  .in1({ S6086, S2832 }),
  .out1({ S39 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4679_ (
  .in1({ S6086, S2843 }),
  .out1({ S40 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4680_ (
  .in1({ S6086, S2854 }),
  .out1({ S41 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4681_ (
  .in1({ S6086, S2865 }),
  .out1({ S42 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4682_ (
  .in1({ S6086, S2876 }),
  .out1({ S43 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4683_ (
  .in1({ S6086, S2887 }),
  .out1({ S44 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4684_ (
  .in1({ S6086, S2898 }),
  .out1({ S45 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4685_ (
  .in1({ S6086, S2909 }),
  .out1({ S46 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4686_ (
  .in1({ S6086, S2920 }),
  .out1({ S47 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4687_ (
  .in1({ S6086, S2931 }),
  .out1({ S48 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4688_ (
  .in1({ S6086, S2942 }),
  .out1({ S49 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4689_ (
  .in1({ S6086, S2953 }),
  .out1({ S50 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4690_ (
  .in1({ new_controller_1133_S_0, new_datapath_databusin_0 }),
  .out1({ S4239 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4691_ (
  .in1({ S6087, new_datapath_instruction_0 }),
  .out1({ S4240 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4692_ (
  .in1({ S4240, S4239 }),
  .out1({ S51 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4693_ (
  .in1({ new_controller_1133_S_0, new_datapath_databusin_1 }),
  .out1({ S4241 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4694_ (
  .in1({ S6087, new_datapath_instruction_1 }),
  .out1({ S4242 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4695_ (
  .in1({ S4242, S4241 }),
  .out1({ S52 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4696_ (
  .in1({ new_controller_1133_S_0, new_datapath_databusin_2 }),
  .out1({ S4243 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4697_ (
  .in1({ S6087, new_datapath_instruction_2 }),
  .out1({ S4244 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4698_ (
  .in1({ S4244, S4243 }),
  .out1({ S53 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4699_ (
  .in1({ new_controller_1133_S_0, new_datapath_databusin_3 }),
  .out1({ S4245 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4700_ (
  .in1({ S6087, new_datapath_instruction_3 }),
  .out1({ S4247 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4701_ (
  .in1({ S4247, S4245 }),
  .out1({ S54 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4702_ (
  .in1({ new_controller_1133_S_0, new_datapath_databusin_4 }),
  .out1({ S4248 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4703_ (
  .in1({ S6087, new_controller_fib_0 }),
  .out1({ S4249 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4704_ (
  .in1({ S4249, S4248 }),
  .out1({ S55 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4705_ (
  .in1({ new_controller_1133_S_0, new_datapath_databusin_5 }),
  .out1({ S4250 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4706_ (
  .in1({ S6087, new_controller_fib_1 }),
  .out1({ S4251 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4707_ (
  .in1({ S4251, S4250 }),
  .out1({ S56 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4708_ (
  .in1({ new_controller_1133_S_0, new_datapath_databusin_6 }),
  .out1({ S4252 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4709_ (
  .in1({ S6087, new_controller_fib_2 }),
  .out1({ S4253 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4710_ (
  .in1({ S4253, S4252 }),
  .out1({ S57 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4711_ (
  .in1({ new_controller_1133_S_0, new_datapath_databusin_7 }),
  .out1({ S4255 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4712_ (
  .in1({ S6087, new_controller_fib_3 }),
  .out1({ S4256 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4713_ (
  .in1({ S4256, S4255 }),
  .out1({ S58 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4714_ (
  .in1({ new_controller_1133_S_0, new_datapath_databusin_8 }),
  .out1({ S4257 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4715_ (
  .in1({ S6087, new_controller_fib_4 }),
  .out1({ S4258 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4716_ (
  .in1({ S4258, S4257 }),
  .out1({ S59 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4717_ (
  .in1({ new_controller_1133_S_0, new_datapath_databusin_9 }),
  .out1({ S4259 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4718_ (
  .in1({ S6087, new_controller_234_B_0 }),
  .out1({ S4260 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4719_ (
  .in1({ S4260, S4259 }),
  .out1({ S60 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4720_ (
  .in1({ new_controller_1133_S_0, new_datapath_databusin_10 }),
  .out1({ S4262 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4721_ (
  .in1({ S6087, new_controller_opcode_2 }),
  .out1({ S4263 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4722_ (
  .in1({ S4263, S4262 }),
  .out1({ S61 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4723_ (
  .in1({ new_controller_1133_S_0, new_datapath_databusin_11 }),
  .out1({ S4264 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4724_ (
  .in1({ S6087, new_controller_opcode_3 }),
  .out1({ S4265 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4725_ (
  .in1({ S4265, S4264 }),
  .out1({ S62 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4726_ (
  .in1({ new_controller_1133_S_0, new_datapath_databusin_12 }),
  .out1({ S4266 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4727_ (
  .in1({ S6087, new_controller_opcode_4 }),
  .out1({ S4267 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4728_ (
  .in1({ S4267, S4266 }),
  .out1({ S63 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4729_ (
  .in1({ new_controller_1133_S_0, new_datapath_databusin_13 }),
  .out1({ S4268 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4730_ (
  .in1({ S6087, new_controller_opcode_5 }),
  .out1({ S4270 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4731_ (
  .in1({ S4270, S4268 }),
  .out1({ S64 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4732_ (
  .in1({ new_controller_1133_S_0, new_datapath_databusin_14 }),
  .out1({ S4271 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4733_ (
  .in1({ S6087, new_controller_opcode_6 }),
  .out1({ S4272 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4734_ (
  .in1({ S4272, S4271 }),
  .out1({ S65 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4735_ (
  .in1({ S172, new_controller_opcode_2 }),
  .out1({ S4273 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4736_ (
  .in1({ S171, S3051 }),
  .out1({ S4274 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4737_ (
  .in1({ S4274, new_controller_407_B_0 }),
  .out1({ S4275 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4738_ (
  .in1({ S4274, S3040 }),
  .out1({ S4276 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4739_ (
  .in1({ S4273, new_controller_234_B_0 }),
  .out1({ S4277 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4740_ (
  .in1({ S4276, S5365 }),
  .out1({ S4279 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4741_ (
  .in1({ S4277, S5354 }),
  .out1({ S4280 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4742_ (
  .in1({ new_datapath_addsubunit_in1_2, S5157 }),
  .out1({ S4281 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4743_ (
  .in1({ S5147, S4067 }),
  .out1({ S4282 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4744_ (
  .in1({ S4282, S3761 }),
  .out1({ S4283 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4745_ (
  .in1({ S4283 }),
  .out1({ S4284 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4746_ (
  .in1({ S4283, S5343 }),
  .out1({ S4285 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4747_ (
  .in1({ S4283, S5354 }),
  .out1({ S4286 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4748_ (
  .in1({ S4284, S4289 }),
  .out1({ S4287 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4749_ (
  .in1({ S4287, S4279 }),
  .out1({ S4288 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4750_ (
  .in1({ S4288, new_controller_fib_2 }),
  .out1({ S4290 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4751_ (
  .in1({ S4290, S4281 }),
  .out1({ S4291 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4752_ (
  .in1({ S4291, S4280 }),
  .out1({ S4292 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4753_ (
  .in1({ S175, S5515 }),
  .out1({ S4293 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4754_ (
  .in1({ S176, S5526 }),
  .out1({ S4294 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4755_ (
  .in1({ S4294, S257 }),
  .out1({ S4295 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4756_ (
  .in1({ S4295, S4292 }),
  .out1({ S4296 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4757_ (
  .in1({ S4296, S5957 }),
  .out1({ S4297 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4758_ (
  .in1({ S4296, new_datapath_addsubunit_in1_2 }),
  .out1({ S4298 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4759_ (
  .in1({ S4298 }),
  .out1({ S4299 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4760_ (
  .in1({ S4296, new_datapath_addsubunit_in1_2 }),
  .out1({ S4301 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4761_ (
  .in1({ S4301, S4299 }),
  .out1({ S4302 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4762_ (
  .in1({ S5907, S5168 }),
  .out1({ S4303 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4763_ (
  .in1({ S4286, new_controller_opcode_3 }),
  .out1({ S4304 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4764_ (
  .in1({ S4276, new_controller_fib_4 }),
  .out1({ S4305 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4765_ (
  .in1({ S4305, S4300 }),
  .out1({ S4306 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4766_ (
  .in1({ S4306 }),
  .out1({ S4307 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4767_ (
  .in1({ S4306, S4303 }),
  .out1({ S4308 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4768_ (
  .in1({ S4308, S4304 }),
  .out1({ S4309 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4769_ (
  .in1({ S4309, S4280 }),
  .out1({ S4310 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4770_ (
  .in1({ S4294, S229 }),
  .out1({ S4312 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4771_ (
  .in1({ S4312, S4310 }),
  .out1({ S4313 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4772_ (
  .in1({ S4313 }),
  .out1({ S4314 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4773_ (
  .in1({ S4314, S5907 }),
  .out1({ S4315 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4774_ (
  .in1({ S4313, new_datapath_addsubunit_in1_7 }),
  .out1({ S4316 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4775_ (
  .in1({ S4313, new_datapath_addsubunit_in1_7 }),
  .out1({ S4317 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4776_ (
  .in1({ S4313, S5907 }),
  .out1({ S4318 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4777_ (
  .in1({ S4314, new_datapath_addsubunit_in1_7 }),
  .out1({ S4319 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4778_ (
  .in1({ S4317, S4315 }),
  .out1({ S4320 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4779_ (
  .in1({ S4320 }),
  .out1({ S4321 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4780_ (
  .in1({ new_datapath_addsubunit_in1_3, S5157 }),
  .out1({ S4323 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4781_ (
  .in1({ S4288, new_controller_fib_3 }),
  .out1({ S4324 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4782_ (
  .in1({ S4324, S4323 }),
  .out1({ S4325 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4783_ (
  .in1({ S4325, S4280 }),
  .out1({ S4326 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4784_ (
  .in1({ S4294, S249 }),
  .out1({ S4327 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4785_ (
  .in1({ S4327, S4326 }),
  .out1({ S4328 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4786_ (
  .in1({ S4328 }),
  .out1({ S4329 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4787_ (
  .in1({ S4329, S5947 }),
  .out1({ S4330 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4788_ (
  .in1({ S4328, new_datapath_addsubunit_in1_3 }),
  .out1({ S4331 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4789_ (
  .in1({ S4328, new_datapath_addsubunit_in1_3 }),
  .out1({ S4332 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4790_ (
  .in1({ S4332 }),
  .out1({ S4334 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4791_ (
  .in1({ S4328, S5947 }),
  .out1({ S4335 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4792_ (
  .in1({ S4329, new_datapath_addsubunit_in1_3 }),
  .out1({ S4336 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4793_ (
  .in1({ S4332, S4330 }),
  .out1({ S4337 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4794_ (
  .in1({ S4334, S4331 }),
  .out1({ S4338 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4795_ (
  .in1({ new_datapath_addsubunit_in1_1, S5157 }),
  .out1({ S4339 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4796_ (
  .in1({ S4288, new_controller_fib_1 }),
  .out1({ S4340 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4797_ (
  .in1({ S4340, S4339 }),
  .out1({ S4341 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4798_ (
  .in1({ S4341, S4280 }),
  .out1({ S4342 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4799_ (
  .in1({ S4294, S265 }),
  .out1({ S4343 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4800_ (
  .in1({ S4343, S4342 }),
  .out1({ S4345 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4801_ (
  .in1({ S4345 }),
  .out1({ S4346 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4802_ (
  .in1({ S4345, S5966 }),
  .out1({ S4347 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4803_ (
  .in1({ S4346, S5966 }),
  .out1({ S4348 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4804_ (
  .in1({ S4345, new_datapath_addsubunit_in1_1 }),
  .out1({ S4349 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4805_ (
  .in1({ S4345, new_datapath_addsubunit_in1_1 }),
  .out1({ S4350 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4806_ (
  .in1({ S4350 }),
  .out1({ S4351 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4807_ (
  .in1({ S4351, S4349 }),
  .out1({ S4352 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4808_ (
  .in1({ S4350, S4348 }),
  .out1({ S4353 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4809_ (
  .in1({ new_datapath_addsubunit_in1_0, S5157 }),
  .out1({ S4354 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4810_ (
  .in1({ S4288, new_controller_fib_0 }),
  .out1({ S4356 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4811_ (
  .in1({ S4356, S4354 }),
  .out1({ S4357 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4812_ (
  .in1({ S4357, S4280 }),
  .out1({ S4358 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4813_ (
  .in1({ S4358 }),
  .out1({ S4359 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4814_ (
  .in1({ S4293, S270 }),
  .out1({ S4360 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4815_ (
  .in1({ S4294, S271 }),
  .out1({ S4361 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4816_ (
  .in1({ S4360, S4359 }),
  .out1({ S4362 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4817_ (
  .in1({ S4361, S4358 }),
  .out1({ S4363 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4818_ (
  .in1({ S4362, new_datapath_addsubunit_in1_0 }),
  .out1({ S4364 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4819_ (
  .in1({ S4364, S4353 }),
  .out1({ S4365 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4820_ (
  .in1({ S5926, S5168 }),
  .out1({ S4367 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4821_ (
  .in1({ S4286, new_controller_234_B_0 }),
  .out1({ S4368 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4822_ (
  .in1({ S4368, S4307 }),
  .out1({ S4369 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4823_ (
  .in1({ S4369, S4367 }),
  .out1({ S4370 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4824_ (
  .in1({ S4370, S4279 }),
  .out1({ S4371 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4825_ (
  .in1({ S4293, S208 }),
  .out1({ S4372 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4826_ (
  .in1({ S4372, S4371 }),
  .out1({ S4373 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4827_ (
  .in1({ S4373 }),
  .out1({ S4374 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4828_ (
  .in1({ S4374, S5926 }),
  .out1({ S4375 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4829_ (
  .in1({ S4373, new_datapath_addsubunit_in1_5 }),
  .out1({ S4376 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4830_ (
  .in1({ S4376, S4375 }),
  .out1({ S4378 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4831_ (
  .in1({ S4378 }),
  .out1({ S4379 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4832_ (
  .in1({ S4363, S5975 }),
  .out1({ S4380 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4833_ (
  .in1({ S4285, new_controller_fib_0 }),
  .out1({ S4381 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4834_ (
  .in1({ S4285, S5157 }),
  .out1({ S4382 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4835_ (
  .in1({ S4382, S3062 }),
  .out1({ S4383 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4836_ (
  .in1({ S4383, S5157 }),
  .out1({ S4384 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4837_ (
  .in1({ S4384, S4381 }),
  .out1({ S4385 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4838_ (
  .in1({ S4385 }),
  .out1({ S4386 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4839_ (
  .in1({ S4385, S4306 }),
  .out1({ S4387 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4840_ (
  .in1({ S4386, S4307 }),
  .out1({ S4389 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4841_ (
  .in1({ S4387, S4279 }),
  .out1({ S4390 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4842_ (
  .in1({ S4389, S4280 }),
  .out1({ S4391 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4843_ (
  .in1({ S4294, new_datapath_multdivunit_1697_B_15 }),
  .out1({ S4392 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4844_ (
  .in1({ S4392 }),
  .out1({ S4393 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4845_ (
  .in1({ S4393, S4390 }),
  .out1({ S4394 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4846_ (
  .in1({ S4394 }),
  .out1({ S4395 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4847_ (
  .in1({ S4394, new_datapath_addsubunit_in1_15 }),
  .out1({ S4396 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4848_ (
  .in1({ S4396 }),
  .out1({ S4397 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4849_ (
  .in1({ S4394, new_datapath_addsubunit_in1_15 }),
  .out1({ S4398 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4850_ (
  .in1({ S4395, S3401 }),
  .out1({ S4400 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4851_ (
  .in1({ S4398, S4397 }),
  .out1({ S4401 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4852_ (
  .in1({ S4294, new_datapath_multdivunit_1697_B_14 }),
  .out1({ S4402 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4853_ (
  .in1({ S4402, S4391 }),
  .out1({ S4403 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4854_ (
  .in1({ S4403 }),
  .out1({ S4404 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4855_ (
  .in1({ S4403, S3390 }),
  .out1({ S4405 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4856_ (
  .in1({ S4404, new_datapath_addsubunit_in1_14 }),
  .out1({ S4406 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4857_ (
  .in1({ S4404, new_datapath_addsubunit_in1_14 }),
  .out1({ S4407 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4858_ (
  .in1({ S4404, S3390 }),
  .out1({ S4408 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4859_ (
  .in1({ S4407, S4405 }),
  .out1({ S4409 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4860_ (
  .in1({ S4409, S4401 }),
  .out1({ S4411 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4861_ (
  .in1({ S4294, new_datapath_multdivunit_1697_B_13 }),
  .out1({ S4412 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4862_ (
  .in1({ S4412, S4391 }),
  .out1({ S4413 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4863_ (
  .in1({ S4413 }),
  .out1({ S4414 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4864_ (
  .in1({ S4413, new_datapath_addsubunit_in1_13 }),
  .out1({ S4415 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4865_ (
  .in1({ S4414, S3379 }),
  .out1({ S4416 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4866_ (
  .in1({ S4416, S4415 }),
  .out1({ S4417 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4867_ (
  .in1({ S4417 }),
  .out1({ S4418 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4868_ (
  .in1({ S4294, new_datapath_multdivunit_1697_B_12 }),
  .out1({ S4419 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4869_ (
  .in1({ S4419 }),
  .out1({ S4420 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4870_ (
  .in1({ S4420, S4390 }),
  .out1({ S4422 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4871_ (
  .in1({ S4419, S4391 }),
  .out1({ S4423 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4872_ (
  .in1({ S4422, S3368 }),
  .out1({ S4424 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4873_ (
  .in1({ S4423, new_datapath_addsubunit_in1_12 }),
  .out1({ S4425 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4874_ (
  .in1({ S4422, new_datapath_addsubunit_in1_12 }),
  .out1({ S4426 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4875_ (
  .in1({ S4425, S4424 }),
  .out1({ S4427 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4876_ (
  .in1({ S4427, S4417 }),
  .out1({ S4428 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4877_ (
  .in1({ S4428 }),
  .out1({ S4429 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4878_ (
  .in1({ S4429, S4411 }),
  .out1({ S4430 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4879_ (
  .in1({ S4294, new_datapath_multdivunit_1697_B_10 }),
  .out1({ S4431 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4880_ (
  .in1({ S4431, S4391 }),
  .out1({ S4433 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4881_ (
  .in1({ S4433, S3346 }),
  .out1({ S4434 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4882_ (
  .in1({ S4433, new_datapath_addsubunit_in1_10 }),
  .out1({ S4435 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4883_ (
  .in1({ S4435 }),
  .out1({ S4436 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4884_ (
  .in1({ S4433, new_datapath_addsubunit_in1_10 }),
  .out1({ S4437 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4885_ (
  .in1({ S4437, S4436 }),
  .out1({ S4438 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4886_ (
  .in1({ S4294, new_datapath_multdivunit_1697_B_8 }),
  .out1({ S4439 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4887_ (
  .in1({ S4439, S4391 }),
  .out1({ S4440 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4888_ (
  .in1({ S4440 }),
  .out1({ S4441 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4889_ (
  .in1({ S4440, new_datapath_addsubunit_in1_8 }),
  .out1({ S4442 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4890_ (
  .in1({ S4442 }),
  .out1({ S4444 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4891_ (
  .in1({ S4440, new_datapath_addsubunit_in1_8 }),
  .out1({ S4445 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4892_ (
  .in1({ S4441, new_datapath_addsubunit_in1_8 }),
  .out1({ S4446 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4893_ (
  .in1({ S4445, S4444 }),
  .out1({ S4447 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4894_ (
  .in1({ S4447 }),
  .out1({ S4448 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4895_ (
  .in1({ S4294, new_datapath_multdivunit_1697_B_9 }),
  .out1({ S4449 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4896_ (
  .in1({ S4449, S4391 }),
  .out1({ S4450 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4897_ (
  .in1({ S4450 }),
  .out1({ S4451 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4898_ (
  .in1({ S4450, S3336 }),
  .out1({ S4452 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4899_ (
  .in1({ S4451, new_datapath_addsubunit_in1_9 }),
  .out1({ S4453 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4900_ (
  .in1({ S4453, S4452 }),
  .out1({ S4455 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4901_ (
  .in1({ S4455 }),
  .out1({ S4456 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4902_ (
  .in1({ S4455, S4448 }),
  .out1({ S4457 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4903_ (
  .in1({ S4294, new_datapath_multdivunit_1697_B_11 }),
  .out1({ S4458 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4904_ (
  .in1({ S4458 }),
  .out1({ S4459 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4905_ (
  .in1({ S4459, S4390 }),
  .out1({ S4460 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4906_ (
  .in1({ S4458, S4391 }),
  .out1({ S4461 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4907_ (
  .in1({ S4460, new_datapath_addsubunit_in1_11 }),
  .out1({ S4462 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4908_ (
  .in1({ S4461, S3357 }),
  .out1({ S4463 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4909_ (
  .in1({ S4460, S3357 }),
  .out1({ S4464 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4910_ (
  .in1({ S4461, new_datapath_addsubunit_in1_11 }),
  .out1({ S4466 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4911_ (
  .in1({ S4466, S4464 }),
  .out1({ S4467 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4912_ (
  .in1({ S5916, S5168 }),
  .out1({ S4468 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4913_ (
  .in1({ S4286, new_controller_opcode_2 }),
  .out1({ S4469 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4914_ (
  .in1({ S4469, S4307 }),
  .out1({ S4470 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4915_ (
  .in1({ S4470, S4468 }),
  .out1({ S4471 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4916_ (
  .in1({ S4471 }),
  .out1({ S4472 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4917_ (
  .in1({ S4472, S4280 }),
  .out1({ S4473 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4918_ (
  .in1({ S4294, S203 }),
  .out1({ S4474 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4919_ (
  .in1({ S4474, S4473 }),
  .out1({ S4475 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4920_ (
  .in1({ S4475 }),
  .out1({ S4477 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4921_ (
  .in1({ S4475, S5916 }),
  .out1({ S4478 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4922_ (
  .in1({ S4477, S5916 }),
  .out1({ S4479 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4923_ (
  .in1({ S4475, new_datapath_addsubunit_in1_6 }),
  .out1({ S4480 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4924_ (
  .in1({ S4475, new_datapath_addsubunit_in1_6 }),
  .out1({ S4481 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4925_ (
  .in1({ S4481, S4479 }),
  .out1({ S4482 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4926_ (
  .in1({ S4482 }),
  .out1({ S4483 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4927_ (
  .in1({ S5936, S5168 }),
  .out1({ S4484 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4928_ (
  .in1({ S4288, new_controller_fib_4 }),
  .out1({ S4485 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4929_ (
  .in1({ S4485 }),
  .out1({ S4486 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4930_ (
  .in1({ S4486, S4484 }),
  .out1({ S4488 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4931_ (
  .in1({ S4488 }),
  .out1({ S4489 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4932_ (
  .in1({ S4488, S4279 }),
  .out1({ S4490 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4933_ (
  .in1({ S4489, S4280 }),
  .out1({ S4491 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4934_ (
  .in1({ S4293, S240 }),
  .out1({ S4492 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4935_ (
  .in1({ S4294, S241 }),
  .out1({ S4493 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4936_ (
  .in1({ S4492, S4490 }),
  .out1({ S4494 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4937_ (
  .in1({ S4493, S4491 }),
  .out1({ S4495 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4938_ (
  .in1({ S4494, S5936 }),
  .out1({ S4496 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4939_ (
  .in1({ S4496 }),
  .out1({ S4497 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4940_ (
  .in1({ S4495, new_datapath_addsubunit_in1_4 }),
  .out1({ S4499 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4941_ (
  .in1({ S4494, new_datapath_addsubunit_in1_4 }),
  .out1({ S4500 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4942_ (
  .in1({ S4499, S4496 }),
  .out1({ S4501 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4943_ (
  .in1({ S4501 }),
  .out1({ S4502 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4944_ (
  .in1({ S4363, new_datapath_addsubunit_in1_0 }),
  .out1({ S4503 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4945_ (
  .in1({ S4380, S4364 }),
  .out1({ S4504 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4946_ (
  .in1({ S4504 }),
  .out1({ S4505 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4947_ (
  .in1({ S4501, S4302 }),
  .out1({ S4506 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4948_ (
  .in1({ S4482, S4320 }),
  .out1({ S4507 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4949_ (
  .in1({ S4506, S4378 }),
  .out1({ S4508 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4950_ (
  .in1({ S4337, S4274 }),
  .out1({ S4510 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4951_ (
  .in1({ S4467, S4438 }),
  .out1({ S4511 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4952_ (
  .in1({ S4511, S4430 }),
  .out1({ S4512 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4953_ (
  .in1({ S4512, S4457 }),
  .out1({ S4513 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4954_ (
  .in1({ S4513, S4504 }),
  .out1({ S4514 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4955_ (
  .in1({ S4514, S4353 }),
  .out1({ S4515 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4956_ (
  .in1({ S4515, S4510 }),
  .out1({ S4516 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4957_ (
  .in1({ S4516, S4508 }),
  .out1({ S4517 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4958_ (
  .in1({ S4517, S4507 }),
  .out1({ S4518 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4959_ (
  .in1({ S4518, S4275 }),
  .out1({ S70 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4960_ (
  .in1({ S4274, new_controller_407_B_2 }),
  .out1({ S4520 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4961_ (
  .in1({ S4365, S4347 }),
  .out1({ S4521 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4962_ (
  .in1({ S4521, S4302 }),
  .out1({ S4522 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4963_ (
  .in1({ S4522, S4297 }),
  .out1({ S4523 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4964_ (
  .in1({ S4523 }),
  .out1({ S4524 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4965_ (
  .in1({ S4523, S4336 }),
  .out1({ S4525 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4966_ (
  .in1({ S4525, S4335 }),
  .out1({ S4526 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4967_ (
  .in1({ S4526 }),
  .out1({ S4527 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4968_ (
  .in1({ S4527, S4502 }),
  .out1({ S4528 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4969_ (
  .in1({ S4528, S4500 }),
  .out1({ S4529 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4970_ (
  .in1({ S4529 }),
  .out1({ S4531 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4971_ (
  .in1({ S4531, S4376 }),
  .out1({ S4532 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4972_ (
  .in1({ S4532, S4375 }),
  .out1({ S4533 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4973_ (
  .in1({ S4533, S4482 }),
  .out1({ S4534 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4974_ (
  .in1({ S4534, S4478 }),
  .out1({ S4535 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4975_ (
  .in1({ S4535 }),
  .out1({ S4536 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4976_ (
  .in1({ S4535, S4319 }),
  .out1({ S4537 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4977_ (
  .in1({ S4537, S4318 }),
  .out1({ S4538 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4978_ (
  .in1({ S4538, S4447 }),
  .out1({ S4539 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4979_ (
  .in1({ S4539 }),
  .out1({ S4540 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4980_ (
  .in1({ S4540, S4446 }),
  .out1({ S4542 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4981_ (
  .in1({ S4542 }),
  .out1({ S4543 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4982_ (
  .in1({ S4543, S4453 }),
  .out1({ S4544 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4983_ (
  .in1({ S4544, S4452 }),
  .out1({ S4545 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4984_ (
  .in1({ S4545, S4438 }),
  .out1({ S4546 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4985_ (
  .in1({ S4546, S4434 }),
  .out1({ S4547 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4986_ (
  .in1({ S4547, S4462 }),
  .out1({ S4548 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4987_ (
  .in1({ S4548, S4463 }),
  .out1({ S4549 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_4988_ (
  .in1({ S4549 }),
  .out1({ S4550 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4989_ (
  .in1({ S4550, S4430 }),
  .out1({ S4551 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4990_ (
  .in1({ S4413, S3379 }),
  .out1({ S4553 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4991_ (
  .in1({ S4414, new_datapath_addsubunit_in1_13 }),
  .out1({ S4554 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4992_ (
  .in1({ S4426, S4417 }),
  .out1({ S4555 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4993_ (
  .in1({ S4555, S4553 }),
  .out1({ S4556 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4994_ (
  .in1({ S4556, S4411 }),
  .out1({ S4557 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4995_ (
  .in1({ S4406, S4396 }),
  .out1({ S4558 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4996_ (
  .in1({ S4558, S4400 }),
  .out1({ S4559 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4997_ (
  .in1({ S4559, S4273 }),
  .out1({ S4560 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_4998_ (
  .in1({ S4560, S4557 }),
  .out1({ S4561 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_4999_ (
  .in1({ S4561, S4551 }),
  .out1({ S4562 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5000_ (
  .in1({ S4562, S4520 }),
  .out1({ S71 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5001_ (
  .in1({ S6091, new_datapath_adr_outreg_0 }),
  .out1({ S4564 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5002_ (
  .in1({ S6090, S5977 }),
  .out1({ S4565 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5003_ (
  .in1({ S4565, S4564 }),
  .out1({ S73 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5004_ (
  .in1({ S6091, new_datapath_adr_outreg_1 }),
  .out1({ S4566 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5005_ (
  .in1({ S6090, S5968 }),
  .out1({ S4567 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5006_ (
  .in1({ S4567, S4566 }),
  .out1({ S74 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5007_ (
  .in1({ S6091, new_datapath_adr_outreg_2 }),
  .out1({ S4568 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5008_ (
  .in1({ S6090, S5959 }),
  .out1({ S4569 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5009_ (
  .in1({ S4569, S4568 }),
  .out1({ S75 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5010_ (
  .in1({ S6091, new_datapath_adr_outreg_3 }),
  .out1({ S4571 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5011_ (
  .in1({ S6090, S5949 }),
  .out1({ S4572 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5012_ (
  .in1({ S4572, S4571 }),
  .out1({ S76 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5013_ (
  .in1({ S6091, new_datapath_adr_outreg_4 }),
  .out1({ S4573 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5014_ (
  .in1({ S6090, S5938 }),
  .out1({ S4574 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5015_ (
  .in1({ S4574, S4573 }),
  .out1({ S77 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5016_ (
  .in1({ S6091, new_datapath_adr_outreg_5 }),
  .out1({ S4575 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5017_ (
  .in1({ S6090, S5928 }),
  .out1({ S4576 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5018_ (
  .in1({ S4576, S4575 }),
  .out1({ S78 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5019_ (
  .in1({ S6091, new_datapath_adr_outreg_6 }),
  .out1({ S4577 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5020_ (
  .in1({ S6090, S5918 }),
  .out1({ S4579 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5021_ (
  .in1({ S4579, S4577 }),
  .out1({ S79 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5022_ (
  .in1({ S6091, new_datapath_adr_outreg_7 }),
  .out1({ S4580 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5023_ (
  .in1({ S6090, S5909 }),
  .out1({ S4581 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5024_ (
  .in1({ S4581, S4580 }),
  .out1({ S80 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5025_ (
  .in1({ S6091, new_datapath_adr_outreg_8 }),
  .out1({ S4582 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5026_ (
  .in1({ S6090, S4975 }),
  .out1({ S4583 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5027_ (
  .in1({ S4583, S4582 }),
  .out1({ S81 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5028_ (
  .in1({ S6091, new_datapath_adr_outreg_9 }),
  .out1({ S4584 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5029_ (
  .in1({ S6090, S4922 }),
  .out1({ S4585 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5030_ (
  .in1({ S4585, S4584 }),
  .out1({ S82 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5031_ (
  .in1({ S6091, new_datapath_adr_outreg_10 }),
  .out1({ S4587 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5032_ (
  .in1({ S6090, S4857 }),
  .out1({ S4588 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5033_ (
  .in1({ S4588, S4587 }),
  .out1({ S83 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5034_ (
  .in1({ S6091, new_datapath_adr_outreg_11 }),
  .out1({ S4589 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5035_ (
  .in1({ S6090, S4804 }),
  .out1({ S4590 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5036_ (
  .in1({ S4590, S4589 }),
  .out1({ S84 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5037_ (
  .in1({ S6091, new_datapath_adr_outreg_12 }),
  .out1({ S4591 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5038_ (
  .in1({ S6090, S4740 }),
  .out1({ S4592 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5039_ (
  .in1({ S4592, S4591 }),
  .out1({ S85 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5040_ (
  .in1({ S6091, new_datapath_adr_outreg_13 }),
  .out1({ S4594 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5041_ (
  .in1({ S6090, S4686 }),
  .out1({ S4595 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5042_ (
  .in1({ S4595, S4594 }),
  .out1({ S86 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5043_ (
  .in1({ S6091, new_datapath_adr_outreg_14 }),
  .out1({ S4596 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5044_ (
  .in1({ S6090, S4621 }),
  .out1({ S4597 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5045_ (
  .in1({ S4597, S4596 }),
  .out1({ S87 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5046_ (
  .in1({ S5136, S4089 }),
  .out1({ S4598 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5047_ (
  .in1({ S4598 }),
  .out1({ S4599 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5048_ (
  .in1({ S5451, S5239 }),
  .out1({ S4600 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5049_ (
  .in1({ S4600 }),
  .out1({ S4601 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5050_ (
  .in1({ S4598, S3870 }),
  .out1({ S4603 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5051_ (
  .in1({ S4600, S5663 }),
  .out1({ S4604 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5052_ (
  .in1({ S4604, S4603 }),
  .out1({ S4605 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5053_ (
  .in1({ S5483, S5311 }),
  .out1({ S4606 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5054_ (
  .in1({ S170, S3947 }),
  .out1({ S4607 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5055_ (
  .in1({ S4607, S4606 }),
  .out1({ S4608 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5056_ (
  .in1({ S4608, S4605 }),
  .out1({ S4609 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5057_ (
  .in1({ S4609, S3761 }),
  .out1({ S4610 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5058_ (
  .in1({ S4166, S3740 }),
  .out1({ S4611 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5059_ (
  .in1({ S4611, S4122 }),
  .out1({ S4612 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5060_ (
  .in1({ S4612, S4610 }),
  .out1({ new_controller_1133_Y })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5061_ (
  .in1({ new_controller_1133_S_0, S6086 }),
  .out1({ S4614 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5062_ (
  .in1({ S4614 }),
  .out1({ new_controller_1423_Y_0 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5063_ (
  .in1({ S4166, S3708 }),
  .out1({ S4615 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5064_ (
  .in1({ S6091, S5611 }),
  .out1({ S4616 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5065_ (
  .in1({ S4616, S6086 }),
  .out1({ S4617 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5066_ (
  .in1({ S4617, S4615 }),
  .out1({ new_controller_1423_Y_1 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5067_ (
  .in1({ S5280, S3620 }),
  .out1({ S4618 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5068_ (
  .in1({ S5271, S3609 }),
  .out1({ S4619 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5069_ (
  .in1({ S4618, S5255 }),
  .out1({ S4620 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5070_ (
  .in1({ S4619, S5262 }),
  .out1({ S4622 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5071_ (
  .in1({ S4620, S3771 }),
  .out1({ S4623 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5072_ (
  .in1({ S4622, S3761 }),
  .out1({ S4624 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5073_ (
  .in1({ S5558, S5280 }),
  .out1({ S4625 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5074_ (
  .in1({ S5568, S5271 }),
  .out1({ S4626 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5075_ (
  .in1({ S4626, S4624 }),
  .out1({ S4627 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5076_ (
  .in1({ S4627, S4505 }),
  .out1({ S4628 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5077_ (
  .in1({ S4600, S3771 }),
  .out1({ S4629 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5078_ (
  .in1({ S4601, S3761 }),
  .out1({ S4630 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5079_ (
  .in1({ S4630, S4503 }),
  .out1({ S4631 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5080_ (
  .in1({ S4598, S3771 }),
  .out1({ S4633 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5081_ (
  .in1({ S4599, S3761 }),
  .out1({ S4634 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5082_ (
  .in1({ S4633, S4357 }),
  .out1({ S4635 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5083_ (
  .in1({ S5975, new_controller_fib_4 }),
  .out1({ S4636 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5084_ (
  .in1({ S4578, S4269 }),
  .out1({ S4637 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5085_ (
  .in1({ S4570, S4278 }),
  .out1({ S4638 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5086_ (
  .in1({ S4637, new_controller_fib_4 }),
  .out1({ S4639 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5087_ (
  .in1({ S4639 }),
  .out1({ S4640 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5088_ (
  .in1({ S4640, S5975 }),
  .out1({ S4641 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5089_ (
  .in1({ S4641 }),
  .out1({ S4642 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5090_ (
  .in1({ S4641, S4637 }),
  .out1({ S4644 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5091_ (
  .in1({ S4644, S4636 }),
  .out1({ S4645 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5092_ (
  .in1({ S241, S5683 }),
  .out1({ S4646 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5093_ (
  .in1({ S5115, new_controller_fib_4 }),
  .out1({ S4647 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5094_ (
  .in1({ S4647, S4646 }),
  .out1({ S4648 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5095_ (
  .in1({ S4648 }),
  .out1({ S4649 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5096_ (
  .in1({ S5632, S3771 }),
  .out1({ S4650 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5097_ (
  .in1({ S5125, S3040 }),
  .out1({ S4651 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5098_ (
  .in1({ S4651, S4650 }),
  .out1({ S4652 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5099_ (
  .in1({ S4652 }),
  .out1({ S4653 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5100_ (
  .in1({ S5653, S3771 }),
  .out1({ S4655 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5101_ (
  .in1({ S5125, new_controller_234_B_0 }),
  .out1({ S4656 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5102_ (
  .in1({ S4656, S4655 }),
  .out1({ S4657 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5103_ (
  .in1({ S4657, S4652 }),
  .out1({ S4658 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5104_ (
  .in1({ S4658 }),
  .out1({ S4659 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5105_ (
  .in1({ S4659, S4648 }),
  .out1({ S4660 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5106_ (
  .in1({ S4658, S4649 }),
  .out1({ S4661 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5107_ (
  .in1({ S4660, new_datapath_shiftunit_1961_A }),
  .out1({ S4662 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5108_ (
  .in1({ S4648, new_datapath_shiftunit_2265_A }),
  .out1({ S4663 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5109_ (
  .in1({ S4663 }),
  .out1({ S4664 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5110_ (
  .in1({ S6215, new_datapath_databusin_0 }),
  .out1({ S4666 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5111_ (
  .in1({ S6086, new_datapath_multdivunit_outmdu1_0 }),
  .out1({ S4667 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5112_ (
  .in1({ S4144, new_datapath_multdivunit_outmdu2_0 }),
  .out1({ S4668 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5113_ (
  .in1({ S170, S4261 }),
  .out1({ S4669 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5114_ (
  .in1({ S4607, S3761 }),
  .out1({ S4670 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5115_ (
  .in1({ S4670, new_datapath_muxmem_in2_0 }),
  .out1({ S4671 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5116_ (
  .in1({ S4668, S4667 }),
  .out1({ S4672 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5117_ (
  .in1({ S4672, S4671 }),
  .out1({ S4673 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5118_ (
  .in1({ S4673, S4666 }),
  .out1({ S4674 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5119_ (
  .in1({ S4674, S4664 }),
  .out1({ S4675 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5120_ (
  .in1({ S4675, S4662 }),
  .out1({ S4677 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5121_ (
  .in1({ S4677, S4645 }),
  .out1({ S4678 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5122_ (
  .in1({ S4678, S4635 }),
  .out1({ S4679 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5123_ (
  .in1({ S4679, S4631 }),
  .out1({ S4680 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5124_ (
  .in1({ S4680, S4628 }),
  .out1({ new_datapath_indatatrf_0 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5125_ (
  .in1({ S4364, S4353 }),
  .out1({ S4681 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5126_ (
  .in1({ S4624, S4365 }),
  .out1({ S4682 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5127_ (
  .in1({ S4682, S4681 }),
  .out1({ S4683 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5128_ (
  .in1({ S4503, S4352 }),
  .out1({ S4684 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5129_ (
  .in1({ S4684 }),
  .out1({ S4685 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5130_ (
  .in1({ S4503, S4352 }),
  .out1({ S4687 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5131_ (
  .in1({ S4687, S4625 }),
  .out1({ S4688 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5132_ (
  .in1({ S4688, S4684 }),
  .out1({ S4689 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5133_ (
  .in1({ S4629, S4348 }),
  .out1({ S4690 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5134_ (
  .in1({ S4644, new_datapath_addsubunit_in1_1 }),
  .out1({ S4691 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5135_ (
  .in1({ S4633, S4341 }),
  .out1({ S4692 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5136_ (
  .in1({ S4641, S5966 }),
  .out1({ S4693 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5137_ (
  .in1({ S4660, new_datapath_shiftunit_1979_A }),
  .out1({ S4694 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5138_ (
  .in1({ S4648, new_datapath_shiftunit_2283_A }),
  .out1({ S4695 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5139_ (
  .in1({ S4144, new_datapath_multdivunit_outmdu2_1 }),
  .out1({ S4696 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5140_ (
  .in1({ S6086, new_datapath_multdivunit_outmdu1_1 }),
  .out1({ S4698 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5141_ (
  .in1({ S4698, S4696 }),
  .out1({ S4699 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5142_ (
  .in1({ S6215, new_datapath_databusin_1 }),
  .out1({ S4700 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5143_ (
  .in1({ S4669, S6110 }),
  .out1({ S4701 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5144_ (
  .in1({ S4701, S4700 }),
  .out1({ S4702 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5145_ (
  .in1({ S4702, S4699 }),
  .out1({ S4703 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5146_ (
  .in1({ S4703, S4695 }),
  .out1({ S4704 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5147_ (
  .in1({ S4704 }),
  .out1({ S4705 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5148_ (
  .in1({ S4705, S4694 }),
  .out1({ S4706 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5149_ (
  .in1({ S4706, S4693 }),
  .out1({ S4707 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5150_ (
  .in1({ S4707, S4692 }),
  .out1({ S4709 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5151_ (
  .in1({ S4641, new_datapath_addsubunit_in1_1 }),
  .out1({ S4710 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5152_ (
  .in1({ S4642, S5966 }),
  .out1({ S4711 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5153_ (
  .in1({ S4709, S4691 }),
  .out1({ S4712 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5154_ (
  .in1({ S4712, S4690 }),
  .out1({ S4713 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5155_ (
  .in1({ S4713, S4689 }),
  .out1({ S4714 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5156_ (
  .in1({ S4714, S4683 }),
  .out1({ new_datapath_indatatrf_1 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5157_ (
  .in1({ S4685, S4349 }),
  .out1({ S4715 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5158_ (
  .in1({ S4715, S4302 }),
  .out1({ S4716 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5159_ (
  .in1({ S4715, S4302 }),
  .out1({ S4717 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5160_ (
  .in1({ S4716, S4625 }),
  .out1({ S4719 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5161_ (
  .in1({ S4719, S4717 }),
  .out1({ S4720 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5162_ (
  .in1({ S4521, S4302 }),
  .out1({ S4721 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5163_ (
  .in1({ S4624, S4522 }),
  .out1({ S4722 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5164_ (
  .in1({ S4722, S4721 }),
  .out1({ S4723 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5165_ (
  .in1({ S4629, S4299 }),
  .out1({ S4724 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5166_ (
  .in1({ S4633, S4291 }),
  .out1({ S4725 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5167_ (
  .in1({ S4661, S3489 }),
  .out1({ S4726 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5168_ (
  .in1({ S4648, new_datapath_shiftunit_2301_A }),
  .out1({ S4727 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5169_ (
  .in1({ S4669, S6124 }),
  .out1({ S4728 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5170_ (
  .in1({ S6086, new_datapath_multdivunit_outmdu1_2 }),
  .out1({ S4730 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5171_ (
  .in1({ S4730, S4728 }),
  .out1({ S4731 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5172_ (
  .in1({ S4144, new_datapath_multdivunit_outmdu2_2 }),
  .out1({ S4732 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5173_ (
  .in1({ S6215, new_datapath_databusin_2 }),
  .out1({ S4733 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5174_ (
  .in1({ S4733, S4732 }),
  .out1({ S4734 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5175_ (
  .in1({ S4734, S4731 }),
  .out1({ S4735 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5176_ (
  .in1({ S4735, S4727 }),
  .out1({ S4736 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5177_ (
  .in1({ S4736, S4726 }),
  .out1({ S4737 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5178_ (
  .in1({ S4737, S4725 }),
  .out1({ S4738 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5179_ (
  .in1({ S4710, S5957 }),
  .out1({ S4739 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5180_ (
  .in1({ S4711, new_datapath_addsubunit_in1_2 }),
  .out1({ S4741 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5181_ (
  .in1({ S4710, S5957 }),
  .out1({ S4742 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5182_ (
  .in1({ S4742, S4637 }),
  .out1({ S4743 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5183_ (
  .in1({ S4743, S4739 }),
  .out1({ S4744 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5184_ (
  .in1({ S4744, S4738 }),
  .out1({ S4745 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5185_ (
  .in1({ S4745, S4724 }),
  .out1({ S4746 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5186_ (
  .in1({ S4746, S4720 }),
  .out1({ S4747 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5187_ (
  .in1({ S4747, S4723 }),
  .out1({ new_datapath_indatatrf_2 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5188_ (
  .in1({ S4523, S4338 }),
  .out1({ S4748 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5189_ (
  .in1({ S4524, S4337 }),
  .out1({ S4749 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5190_ (
  .in1({ S4749, S4748 }),
  .out1({ S4751 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5191_ (
  .in1({ S4751, S4624 }),
  .out1({ S4752 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5192_ (
  .in1({ S4716, S4298 }),
  .out1({ S4753 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5193_ (
  .in1({ S4753 }),
  .out1({ S4754 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5194_ (
  .in1({ S4753, S4338 }),
  .out1({ S4755 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5195_ (
  .in1({ S4754, S4337 }),
  .out1({ S4756 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5196_ (
  .in1({ S4756, S4755 }),
  .out1({ S4757 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5197_ (
  .in1({ S4757, S4625 }),
  .out1({ S4758 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5198_ (
  .in1({ S4742, new_datapath_addsubunit_in1_3 }),
  .out1({ S4759 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5199_ (
  .in1({ S4742, new_datapath_addsubunit_in1_3 }),
  .out1({ S4760 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5200_ (
  .in1({ S4741, S5947 }),
  .out1({ S4762 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5201_ (
  .in1({ S4760, S4638 }),
  .out1({ S4763 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5202_ (
  .in1({ S4763, S4759 }),
  .out1({ S4764 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5203_ (
  .in1({ S4630, S4331 }),
  .out1({ S4765 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5204_ (
  .in1({ S4633, S4325 }),
  .out1({ S4766 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5205_ (
  .in1({ S4661, S3500 }),
  .out1({ S4767 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5206_ (
  .in1({ S4648, new_datapath_shiftunit_2319_A }),
  .out1({ S4768 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5207_ (
  .in1({ S4669, S6140 }),
  .out1({ S4769 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5208_ (
  .in1({ S6215, new_datapath_databusin_3 }),
  .out1({ S4770 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5209_ (
  .in1({ S4770, S4769 }),
  .out1({ S4771 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5210_ (
  .in1({ S6086, new_datapath_multdivunit_outmdu1_3 }),
  .out1({ S4773 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5211_ (
  .in1({ S4144, new_datapath_multdivunit_outmdu2_3 }),
  .out1({ S4774 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5212_ (
  .in1({ S4774, S4773 }),
  .out1({ S4775 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5213_ (
  .in1({ S4775, S4771 }),
  .out1({ S4776 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5214_ (
  .in1({ S4776, S4768 }),
  .out1({ S4777 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5215_ (
  .in1({ S4777, S4767 }),
  .out1({ S4778 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5216_ (
  .in1({ S4778, S4766 }),
  .out1({ S4779 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5217_ (
  .in1({ S4779, S4765 }),
  .out1({ S4780 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5218_ (
  .in1({ S4780, S4764 }),
  .out1({ S4781 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5219_ (
  .in1({ S4781, S4752 }),
  .out1({ S4782 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5220_ (
  .in1({ S4782, S4758 }),
  .out1({ new_datapath_indatatrf_3 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5221_ (
  .in1({ S4526, S4501 }),
  .out1({ S4784 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5222_ (
  .in1({ S4784, S4528 }),
  .out1({ S4785 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5223_ (
  .in1({ S4785, S4624 }),
  .out1({ S4786 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5224_ (
  .in1({ S4753, S4334 }),
  .out1({ S4787 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5225_ (
  .in1({ S4787, S4331 }),
  .out1({ S4788 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5226_ (
  .in1({ S4788, S4501 }),
  .out1({ S4789 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5227_ (
  .in1({ S4788, S4501 }),
  .out1({ S4790 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5228_ (
  .in1({ S4789, S4626 }),
  .out1({ S4791 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5229_ (
  .in1({ S4791, S4790 }),
  .out1({ S4792 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5230_ (
  .in1({ S4760, S5936 }),
  .out1({ S4794 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5231_ (
  .in1({ S4762, new_datapath_addsubunit_in1_4 }),
  .out1({ S4795 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5232_ (
  .in1({ S4760, S5936 }),
  .out1({ S4796 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5233_ (
  .in1({ S4796, S4637 }),
  .out1({ S4797 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5234_ (
  .in1({ S4797, S4794 }),
  .out1({ S4798 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5235_ (
  .in1({ S4629, S4496 }),
  .out1({ S4799 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5236_ (
  .in1({ S4634, S4488 }),
  .out1({ S4800 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5237_ (
  .in1({ S4660, new_datapath_shiftunit_2033_A }),
  .out1({ S4801 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5238_ (
  .in1({ S4648, new_datapath_shiftunit_2337_A }),
  .out1({ S4802 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5239_ (
  .in1({ S6215, new_datapath_databusin_4 }),
  .out1({ S4803 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5240_ (
  .in1({ S6086, new_datapath_multdivunit_outmdu1_4 }),
  .out1({ S4805 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5241_ (
  .in1({ S4144, new_datapath_multdivunit_outmdu2_4 }),
  .out1({ S4806 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5242_ (
  .in1({ S4670, S6153 }),
  .out1({ S4807 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5243_ (
  .in1({ S4806, S4805 }),
  .out1({ S4808 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5244_ (
  .in1({ S4808, S4807 }),
  .out1({ S4809 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5245_ (
  .in1({ S4809, S4802 }),
  .out1({ S4810 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5246_ (
  .in1({ S4810 }),
  .out1({ S4811 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5247_ (
  .in1({ S4811, S4801 }),
  .out1({ S4812 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5248_ (
  .in1({ S4812, S4800 }),
  .out1({ S4813 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5249_ (
  .in1({ S4813, S4799 }),
  .out1({ S4814 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5250_ (
  .in1({ S4814, S4798 }),
  .out1({ S4816 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5251_ (
  .in1({ S4816, S4803 }),
  .out1({ S4817 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5252_ (
  .in1({ S4817, S4786 }),
  .out1({ S4818 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5253_ (
  .in1({ S4818, S4792 }),
  .out1({ new_datapath_indatatrf_4 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5254_ (
  .in1({ S4529, S4378 }),
  .out1({ S4819 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5255_ (
  .in1({ S4529, S4378 }),
  .out1({ S4820 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5256_ (
  .in1({ S4820, S4623 }),
  .out1({ S4821 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5257_ (
  .in1({ S4821, S4819 }),
  .out1({ S4822 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5258_ (
  .in1({ S4790, S4497 }),
  .out1({ S4823 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5259_ (
  .in1({ S4823, S4379 }),
  .out1({ S4824 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5260_ (
  .in1({ S4824 }),
  .out1({ S4826 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5261_ (
  .in1({ S4823, S4379 }),
  .out1({ S4827 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5262_ (
  .in1({ S4824, S4625 }),
  .out1({ S4828 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5263_ (
  .in1({ S4828, S4827 }),
  .out1({ S4829 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5264_ (
  .in1({ S4373, S5926 }),
  .out1({ S4830 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5265_ (
  .in1({ S4830, S4629 }),
  .out1({ S4831 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5266_ (
  .in1({ S4634, S4370 }),
  .out1({ S4832 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5267_ (
  .in1({ S4660, new_datapath_shiftunit_2051_A }),
  .out1({ S4833 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5268_ (
  .in1({ S4648, new_datapath_shiftunit_2355_A }),
  .out1({ S4834 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5269_ (
  .in1({ S4834 }),
  .out1({ S4835 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5270_ (
  .in1({ S4670, S6167 }),
  .out1({ S4837 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5271_ (
  .in1({ S4144, new_datapath_multdivunit_outmdu2_5 }),
  .out1({ S4838 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5272_ (
  .in1({ S6215, new_datapath_databusin_5 }),
  .out1({ S4839 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5273_ (
  .in1({ S6086, new_datapath_multdivunit_outmdu1_5 }),
  .out1({ S4840 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5274_ (
  .in1({ S4840, S4838 }),
  .out1({ S4841 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5275_ (
  .in1({ S4841, S4837 }),
  .out1({ S4842 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5276_ (
  .in1({ S4842, S4839 }),
  .out1({ S4843 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5277_ (
  .in1({ S4843, S4835 }),
  .out1({ S4844 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5278_ (
  .in1({ S4844, S4833 }),
  .out1({ S4845 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5279_ (
  .in1({ S4845, S4832 }),
  .out1({ S4846 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5280_ (
  .in1({ S4846, S4831 }),
  .out1({ S4848 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5281_ (
  .in1({ S4796, new_datapath_addsubunit_in1_5 }),
  .out1({ S4849 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5282_ (
  .in1({ S4795, S5926 }),
  .out1({ S4850 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5283_ (
  .in1({ S4850 }),
  .out1({ S4851 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5284_ (
  .in1({ S4849, S4637 }),
  .out1({ S4852 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5285_ (
  .in1({ S4852, S4851 }),
  .out1({ S4853 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5286_ (
  .in1({ S4853, S4822 }),
  .out1({ S4854 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5287_ (
  .in1({ S4848, S4829 }),
  .out1({ S4855 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5288_ (
  .in1({ S4855, S4854 }),
  .out1({ new_datapath_indatatrf_5 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5289_ (
  .in1({ S4533, S4482 }),
  .out1({ S4856 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5290_ (
  .in1({ S4856, S4623 }),
  .out1({ S4858 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5291_ (
  .in1({ S4858, S4534 }),
  .out1({ S4859 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5292_ (
  .in1({ S4830, S4826 }),
  .out1({ S4860 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5293_ (
  .in1({ S4860, S4483 }),
  .out1({ S4861 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5294_ (
  .in1({ S4860, S4483 }),
  .out1({ S4862 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5295_ (
  .in1({ S4862 }),
  .out1({ S4863 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5296_ (
  .in1({ S4862, S4626 }),
  .out1({ S4864 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5297_ (
  .in1({ S4864, S4861 }),
  .out1({ S4865 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5298_ (
  .in1({ S4850, new_datapath_addsubunit_in1_6 }),
  .out1({ S4866 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5299_ (
  .in1({ S4850, new_datapath_addsubunit_in1_6 }),
  .out1({ S4867 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5300_ (
  .in1({ S4867, S4638 }),
  .out1({ S4869 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5301_ (
  .in1({ S4869, S4866 }),
  .out1({ S4870 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5302_ (
  .in1({ S4630, S4480 }),
  .out1({ S4871 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5303_ (
  .in1({ S4633, S4472 }),
  .out1({ S4872 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5304_ (
  .in1({ S4661, S3511 }),
  .out1({ S4873 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5305_ (
  .in1({ S4648, new_datapath_shiftunit_2373_A }),
  .out1({ S4874 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5306_ (
  .in1({ S4670, S6179 }),
  .out1({ S4875 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5307_ (
  .in1({ S6086, new_datapath_multdivunit_outmdu1_6 }),
  .out1({ S4876 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5308_ (
  .in1({ S6215, new_datapath_databusin_6 }),
  .out1({ S4877 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5309_ (
  .in1({ S4144, new_datapath_multdivunit_outmdu2_6 }),
  .out1({ S4878 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5310_ (
  .in1({ S4878, S4877 }),
  .out1({ S4880 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5311_ (
  .in1({ S4880 }),
  .out1({ S4881 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5312_ (
  .in1({ S4881, S4876 }),
  .out1({ S4882 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5313_ (
  .in1({ S4882, S4875 }),
  .out1({ S4883 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5314_ (
  .in1({ S4883, S4874 }),
  .out1({ S4884 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5315_ (
  .in1({ S4884, S4873 }),
  .out1({ S4885 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5316_ (
  .in1({ S4885, S4872 }),
  .out1({ S4886 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5317_ (
  .in1({ S4886, S4871 }),
  .out1({ S4887 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5318_ (
  .in1({ S4887, S4870 }),
  .out1({ S4888 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5319_ (
  .in1({ S4888, S4859 }),
  .out1({ S4889 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5320_ (
  .in1({ S4889, S4865 }),
  .out1({ new_datapath_indatatrf_6 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5321_ (
  .in1({ S4535, S4321 }),
  .out1({ S4891 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5322_ (
  .in1({ S4536, S4320 }),
  .out1({ S4892 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5323_ (
  .in1({ S4892, S4891 }),
  .out1({ S4893 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5324_ (
  .in1({ S4893, S4624 }),
  .out1({ S4894 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5325_ (
  .in1({ S4863, S4480 }),
  .out1({ S4895 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5326_ (
  .in1({ S4895, S4320 }),
  .out1({ S4896 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5327_ (
  .in1({ S4895, S4320 }),
  .out1({ S4897 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5328_ (
  .in1({ S4897 }),
  .out1({ S4898 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5329_ (
  .in1({ S4898, S4896 }),
  .out1({ S4899 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5330_ (
  .in1({ S4899, S4625 }),
  .out1({ S4901 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5331_ (
  .in1({ S4630, S4316 }),
  .out1({ S4902 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5332_ (
  .in1({ S4633, S4309 }),
  .out1({ S4903 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5333_ (
  .in1({ S4661, S3522 }),
  .out1({ S4904 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5334_ (
  .in1({ S4648, new_datapath_shiftunit_2391_A }),
  .out1({ S4905 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5335_ (
  .in1({ S4905 }),
  .out1({ S4906 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5336_ (
  .in1({ S4670, S6193 }),
  .out1({ S4907 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5337_ (
  .in1({ S6086, new_datapath_multdivunit_outmdu1_7 }),
  .out1({ S4908 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5338_ (
  .in1({ S6215, new_datapath_databusin_7 }),
  .out1({ S4909 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5339_ (
  .in1({ S4144, new_datapath_multdivunit_outmdu2_7 }),
  .out1({ S4910 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5340_ (
  .in1({ S4910, S4908 }),
  .out1({ S4912 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5341_ (
  .in1({ S4912, S4907 }),
  .out1({ S4913 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5342_ (
  .in1({ S4913, S4909 }),
  .out1({ S4914 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5343_ (
  .in1({ S4914, S4906 }),
  .out1({ S4915 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5344_ (
  .in1({ S4867, S5907 }),
  .out1({ S4916 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5345_ (
  .in1({ S4867, S5907 }),
  .out1({ S4917 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5346_ (
  .in1({ S4917, S4637 }),
  .out1({ S4918 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5347_ (
  .in1({ S4918, S4916 }),
  .out1({ S4919 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5348_ (
  .in1({ S4915, S4903 }),
  .out1({ S4920 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5349_ (
  .in1({ S4920, S4902 }),
  .out1({ S4921 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5350_ (
  .in1({ S4919, S4904 }),
  .out1({ S4923 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5351_ (
  .in1({ S4923, S4921 }),
  .out1({ S4924 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5352_ (
  .in1({ S4924, S4894 }),
  .out1({ S4925 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5353_ (
  .in1({ S4925, S4901 }),
  .out1({ new_datapath_indatatrf_7 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5354_ (
  .in1({ S4538, S4447 }),
  .out1({ S4926 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5355_ (
  .in1({ S4926, S4623 }),
  .out1({ S4927 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5356_ (
  .in1({ S4927, S4539 }),
  .out1({ S4928 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5357_ (
  .in1({ S4895, S4315 }),
  .out1({ S4929 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5358_ (
  .in1({ S4929, S4317 }),
  .out1({ S4930 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5359_ (
  .in1({ S4930, S4447 }),
  .out1({ S4931 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5360_ (
  .in1({ S4930, S4447 }),
  .out1({ S4933 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5361_ (
  .in1({ S4933, S4626 }),
  .out1({ S4934 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5362_ (
  .in1({ S4934, S4931 }),
  .out1({ S4935 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5363_ (
  .in1({ S4917, new_datapath_addsubunit_in1_8 }),
  .out1({ S4936 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5364_ (
  .in1({ S4917, new_datapath_addsubunit_in1_8 }),
  .out1({ S4937 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5365_ (
  .in1({ S4937, S4638 }),
  .out1({ S4938 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5366_ (
  .in1({ S4938, S4936 }),
  .out1({ S4939 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5367_ (
  .in1({ S4661, S3533 }),
  .out1({ S4940 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5368_ (
  .in1({ S4648, new_datapath_shiftunit_2409_A }),
  .out1({ S4941 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5369_ (
  .in1({ S4629, S4444 }),
  .out1({ S4942 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5370_ (
  .in1({ S4633, S4389 }),
  .out1({ S4944 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5371_ (
  .in1({ S4670, S6205 }),
  .out1({ S4945 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5372_ (
  .in1({ S6086, new_datapath_multdivunit_outmdu1_8 }),
  .out1({ S4946 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5373_ (
  .in1({ S6215, new_datapath_databusin_8 }),
  .out1({ S4947 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5374_ (
  .in1({ S4144, new_datapath_multdivunit_outmdu2_8 }),
  .out1({ S4948 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5375_ (
  .in1({ S4947, S4944 }),
  .out1({ S4949 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5376_ (
  .in1({ S4948, S4946 }),
  .out1({ S4950 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5377_ (
  .in1({ S4950, S4945 }),
  .out1({ S4951 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5378_ (
  .in1({ S4951, S4942 }),
  .out1({ S4952 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5379_ (
  .in1({ S4952, S4949 }),
  .out1({ S4953 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5380_ (
  .in1({ S4953, S4941 }),
  .out1({ S4955 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5381_ (
  .in1({ S4955, S4940 }),
  .out1({ S4956 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5382_ (
  .in1({ S4956, S4939 }),
  .out1({ S4957 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5383_ (
  .in1({ S4957, S4928 }),
  .out1({ S4958 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5384_ (
  .in1({ S4958, S4935 }),
  .out1({ new_datapath_indatatrf_8 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5385_ (
  .in1({ S4542, S4455 }),
  .out1({ S4959 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5386_ (
  .in1({ S4543, S4456 }),
  .out1({ S4960 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5387_ (
  .in1({ S4960, S4959 }),
  .out1({ S4961 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5388_ (
  .in1({ S4961, S4623 }),
  .out1({ S4962 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5389_ (
  .in1({ S4931, S4442 }),
  .out1({ S4963 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5390_ (
  .in1({ S4963, S4456 }),
  .out1({ S4965 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5391_ (
  .in1({ S4963, S4456 }),
  .out1({ S4966 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5392_ (
  .in1({ S4966, S4625 }),
  .out1({ S4967 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5393_ (
  .in1({ S4967, S4965 }),
  .out1({ S4968 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5394_ (
  .in1({ S4937, S3336 }),
  .out1({ S4969 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5395_ (
  .in1({ S4937, S3336 }),
  .out1({ S4970 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5396_ (
  .in1({ S4970, S4637 }),
  .out1({ S4971 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5397_ (
  .in1({ S4971, S4969 }),
  .out1({ S4972 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5398_ (
  .in1({ S4661, S3544 }),
  .out1({ S4973 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5399_ (
  .in1({ S4648, new_datapath_shiftunit_2427_A }),
  .out1({ S4974 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5400_ (
  .in1({ S4450, new_datapath_addsubunit_in1_9 }),
  .out1({ S4976 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5401_ (
  .in1({ S4976, S4630 }),
  .out1({ S4977 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5402_ (
  .in1({ S4285, new_controller_fib_1 }),
  .out1({ S4978 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5403_ (
  .in1({ S4978, S4384 }),
  .out1({ S4979 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5404_ (
  .in1({ S4979, S4306 }),
  .out1({ S4980 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5405_ (
  .in1({ S4980, S4634 }),
  .out1({ S4981 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5406_ (
  .in1({ S4669, S93 }),
  .out1({ S4982 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5407_ (
  .in1({ S6086, new_datapath_multdivunit_outmdu1_9 }),
  .out1({ S4983 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5408_ (
  .in1({ S6215, new_datapath_databusin_9 }),
  .out1({ S4984 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5409_ (
  .in1({ S4144, new_datapath_multdivunit_outmdu2_9 }),
  .out1({ S4985 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5410_ (
  .in1({ S4985, S4983 }),
  .out1({ S4987 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5411_ (
  .in1({ S4987, S4981 }),
  .out1({ S4988 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5412_ (
  .in1({ S4988, S4982 }),
  .out1({ S4989 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5413_ (
  .in1({ S4989, S4977 }),
  .out1({ S4990 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5414_ (
  .in1({ S4990, S4984 }),
  .out1({ S4991 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5415_ (
  .in1({ S4991, S4973 }),
  .out1({ S4992 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5416_ (
  .in1({ S4992, S4974 }),
  .out1({ S4993 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5417_ (
  .in1({ S4993, S4972 }),
  .out1({ S4994 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5418_ (
  .in1({ S4994 }),
  .out1({ S4995 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5419_ (
  .in1({ S4995, S4968 }),
  .out1({ S4996 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5420_ (
  .in1({ S4996, S4962 }),
  .out1({ new_datapath_indatatrf_9 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5421_ (
  .in1({ S4545, S4438 }),
  .out1({ S4998 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5422_ (
  .in1({ S4624, S4546 }),
  .out1({ S4999 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5423_ (
  .in1({ S4999, S4998 }),
  .out1({ S5000 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5424_ (
  .in1({ S4976, S4966 }),
  .out1({ S5001 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5425_ (
  .in1({ S5001, S4438 }),
  .out1({ S5002 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5426_ (
  .in1({ S5001, S4438 }),
  .out1({ S5003 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5427_ (
  .in1({ S5003, S4625 }),
  .out1({ S5004 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5428_ (
  .in1({ S5004, S5002 }),
  .out1({ S5005 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5429_ (
  .in1({ S4970, new_datapath_addsubunit_in1_10 }),
  .out1({ S5006 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5430_ (
  .in1({ S4970, new_datapath_addsubunit_in1_10 }),
  .out1({ S5008 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5431_ (
  .in1({ S5008 }),
  .out1({ S5009 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5432_ (
  .in1({ S5008, S4638 }),
  .out1({ S5010 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5433_ (
  .in1({ S5010, S5006 }),
  .out1({ S5011 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5434_ (
  .in1({ S4661, S3554 }),
  .out1({ S5012 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5435_ (
  .in1({ S4648, new_datapath_shiftunit_2445_A }),
  .out1({ S5013 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5436_ (
  .in1({ S4630, S4435 }),
  .out1({ S5014 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5437_ (
  .in1({ S4669, S107 }),
  .out1({ S5015 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5438_ (
  .in1({ S4285, new_controller_fib_2 }),
  .out1({ S5016 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5439_ (
  .in1({ S5016, S4384 }),
  .out1({ S5017 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5440_ (
  .in1({ S5017, S4306 }),
  .out1({ S5019 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5441_ (
  .in1({ S5019, S4634 }),
  .out1({ S5020 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5442_ (
  .in1({ S4144, new_datapath_multdivunit_outmdu2_10 }),
  .out1({ S5021 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5443_ (
  .in1({ S6086, new_datapath_multdivunit_outmdu1_10 }),
  .out1({ S5022 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5444_ (
  .in1({ S6215, new_datapath_databusin_10 }),
  .out1({ S5023 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5445_ (
  .in1({ S5023, S5022 }),
  .out1({ S5024 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5446_ (
  .in1({ S5024 }),
  .out1({ S5025 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5447_ (
  .in1({ S5025, S5021 }),
  .out1({ S5026 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5448_ (
  .in1({ S5026, S5020 }),
  .out1({ S5027 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5449_ (
  .in1({ S5027, S5015 }),
  .out1({ S5028 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5450_ (
  .in1({ S5028, S5014 }),
  .out1({ S5030 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5451_ (
  .in1({ S5030, S5013 }),
  .out1({ S5031 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5452_ (
  .in1({ S5031, S5012 }),
  .out1({ S5032 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5453_ (
  .in1({ S5032, S5011 }),
  .out1({ S5033 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5454_ (
  .in1({ S5033, S5005 }),
  .out1({ S5034 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5455_ (
  .in1({ S5034, S5000 }),
  .out1({ new_datapath_indatatrf_10 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5456_ (
  .in1({ S4547, S4467 }),
  .out1({ S5035 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5457_ (
  .in1({ S4547, S4467 }),
  .out1({ S5036 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5458_ (
  .in1({ S5036 }),
  .out1({ S5037 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5459_ (
  .in1({ S5037, S5035 }),
  .out1({ S5038 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5460_ (
  .in1({ S5038, S4624 }),
  .out1({ S5040 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5461_ (
  .in1({ S5003, S4435 }),
  .out1({ S5041 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5462_ (
  .in1({ S5041, S4467 }),
  .out1({ S5042 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5463_ (
  .in1({ S5042 }),
  .out1({ S5043 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5464_ (
  .in1({ S5041, S4467 }),
  .out1({ S5044 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5465_ (
  .in1({ S5044, S5043 }),
  .out1({ S5045 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5466_ (
  .in1({ S5045, S4626 }),
  .out1({ S5046 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5467_ (
  .in1({ S4661, S3565 }),
  .out1({ S5047 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5468_ (
  .in1({ S4648, new_datapath_shiftunit_2463_A }),
  .out1({ S5048 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5469_ (
  .in1({ S4629, S4464 }),
  .out1({ S5049 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5470_ (
  .in1({ S4670, S122 }),
  .out1({ S5051 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5471_ (
  .in1({ S4285, new_controller_fib_3 }),
  .out1({ S5052 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5472_ (
  .in1({ S5052, S4384 }),
  .out1({ S5053 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5473_ (
  .in1({ S5053, S4306 }),
  .out1({ S5054 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5474_ (
  .in1({ S5054, S4634 }),
  .out1({ S5055 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5475_ (
  .in1({ S4144, new_datapath_multdivunit_outmdu2_11 }),
  .out1({ S5056 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5476_ (
  .in1({ S6215, new_datapath_databusin_11 }),
  .out1({ S5057 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5477_ (
  .in1({ S5057, S5056 }),
  .out1({ S5058 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5478_ (
  .in1({ S6086, new_datapath_multdivunit_outmdu1_11 }),
  .out1({ S5059 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5479_ (
  .in1({ S5055, S5051 }),
  .out1({ S5060 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5480_ (
  .in1({ S5059, S5049 }),
  .out1({ S5062 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5481_ (
  .in1({ S5062, S5058 }),
  .out1({ S5063 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5482_ (
  .in1({ S5063, S5048 }),
  .out1({ S5064 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5483_ (
  .in1({ S5064, S5047 }),
  .out1({ S5065 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5484_ (
  .in1({ S5065, S5060 }),
  .out1({ S5066 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5485_ (
  .in1({ S5009, new_datapath_addsubunit_in1_11 }),
  .out1({ S5067 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5486_ (
  .in1({ S5008, S3357 }),
  .out1({ S5068 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5487_ (
  .in1({ S5068, S5067 }),
  .out1({ S5069 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5488_ (
  .in1({ S5069, S4638 }),
  .out1({ S5070 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5489_ (
  .in1({ S5066, S5040 }),
  .out1({ S5071 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5490_ (
  .in1({ S5070, S5046 }),
  .out1({ S5073 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5491_ (
  .in1({ S5073, S5071 }),
  .out1({ new_datapath_indatatrf_11 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5492_ (
  .in1({ S4549, S4427 }),
  .out1({ S5074 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5493_ (
  .in1({ S4549, S4427 }),
  .out1({ S5075 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5494_ (
  .in1({ S5075 }),
  .out1({ S5076 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5495_ (
  .in1({ S5075, S4624 }),
  .out1({ S5077 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5496_ (
  .in1({ S5077, S5074 }),
  .out1({ S5078 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5497_ (
  .in1({ S5041, S4464 }),
  .out1({ S5079 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5498_ (
  .in1({ S5079, S4466 }),
  .out1({ S5080 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5499_ (
  .in1({ S5080, S4427 }),
  .out1({ S5081 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5500_ (
  .in1({ S5080, S4427 }),
  .out1({ S5083 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5501_ (
  .in1({ S5083 }),
  .out1({ S5084 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5502_ (
  .in1({ S5083, S4625 }),
  .out1({ S5085 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5503_ (
  .in1({ S5085, S5081 }),
  .out1({ S5086 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5504_ (
  .in1({ S5068, new_datapath_addsubunit_in1_12 }),
  .out1({ S5087 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5505_ (
  .in1({ S5068, new_datapath_addsubunit_in1_12 }),
  .out1({ S5088 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5506_ (
  .in1({ S5088 }),
  .out1({ S5089 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5507_ (
  .in1({ S5088, S4638 }),
  .out1({ S5090 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5508_ (
  .in1({ S5090, S5087 }),
  .out1({ S5091 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5509_ (
  .in1({ S4661, S3576 }),
  .out1({ S5092 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5510_ (
  .in1({ S4648, new_datapath_shiftunit_2481_A }),
  .out1({ S5094 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5511_ (
  .in1({ S4670, S134 }),
  .out1({ S5095 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5512_ (
  .in1({ S4629, S4424 }),
  .out1({ S5096 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5513_ (
  .in1({ S4285, new_controller_fib_4 }),
  .out1({ S5097 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5514_ (
  .in1({ S5097, S4384 }),
  .out1({ S5098 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5515_ (
  .in1({ S5098, S4306 }),
  .out1({ S5099 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5516_ (
  .in1({ S5099, S4634 }),
  .out1({ S5100 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5517_ (
  .in1({ S4144, new_datapath_multdivunit_outmdu2_12 }),
  .out1({ S5101 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5518_ (
  .in1({ S6215, new_datapath_databusin_12 }),
  .out1({ S5102 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5519_ (
  .in1({ S6086, new_datapath_multdivunit_outmdu1_12 }),
  .out1({ S5103 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5520_ (
  .in1({ S5103, S5102 }),
  .out1({ S5105 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5521_ (
  .in1({ S5105 }),
  .out1({ S5106 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5522_ (
  .in1({ S5106, S5101 }),
  .out1({ S5107 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5523_ (
  .in1({ S5107, S5100 }),
  .out1({ S5108 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5524_ (
  .in1({ S5108, S5096 }),
  .out1({ S5109 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5525_ (
  .in1({ S5109, S5095 }),
  .out1({ S5110 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5526_ (
  .in1({ S5110, S5094 }),
  .out1({ S5111 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5527_ (
  .in1({ S5111, S5092 }),
  .out1({ S5112 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5528_ (
  .in1({ S5112, S5091 }),
  .out1({ S5113 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5529_ (
  .in1({ S5113, S5086 }),
  .out1({ S5114 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5530_ (
  .in1({ S5114, S5078 }),
  .out1({ new_datapath_indatatrf_12 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5531_ (
  .in1({ S5076, S4426 }),
  .out1({ S5116 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5532_ (
  .in1({ S5116, S4418 }),
  .out1({ S5117 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5533_ (
  .in1({ S5116, S4418 }),
  .out1({ S5118 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5534_ (
  .in1({ S5118, S4624 }),
  .out1({ S5119 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5535_ (
  .in1({ S5119, S5117 }),
  .out1({ S5120 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5536_ (
  .in1({ S5084, S4424 }),
  .out1({ S5121 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5537_ (
  .in1({ S5121, S4417 }),
  .out1({ S5122 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5538_ (
  .in1({ S5121, S4417 }),
  .out1({ S5123 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5539_ (
  .in1({ S5123 }),
  .out1({ S5124 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5540_ (
  .in1({ S5124, S5122 }),
  .out1({ S5126 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5541_ (
  .in1({ S5126, S4626 }),
  .out1({ S5127 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5542_ (
  .in1({ S5088, S3379 }),
  .out1({ S5128 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5543_ (
  .in1({ S5089, new_datapath_addsubunit_in1_13 }),
  .out1({ S5129 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5544_ (
  .in1({ S5129 }),
  .out1({ S5130 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5545_ (
  .in1({ S5129, S5128 }),
  .out1({ S5131 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5546_ (
  .in1({ S5131, S4637 }),
  .out1({ S5132 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5547_ (
  .in1({ S4660, new_datapath_shiftunit_2195_A }),
  .out1({ S5133 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5548_ (
  .in1({ S4648, new_datapath_shiftunit_2499_A }),
  .out1({ S5134 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5549_ (
  .in1({ S4670, S148 }),
  .out1({ S5135 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5550_ (
  .in1({ S4629, S4416 }),
  .out1({ S5137 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5551_ (
  .in1({ S4285, new_controller_234_B_0 }),
  .out1({ S5138 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5552_ (
  .in1({ S5138, S4384 }),
  .out1({ S5139 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5553_ (
  .in1({ S5139, S4306 }),
  .out1({ S5140 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5554_ (
  .in1({ S5140, S4634 }),
  .out1({ S5141 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5555_ (
  .in1({ S4144, new_datapath_multdivunit_outmdu2_13 }),
  .out1({ S5142 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5556_ (
  .in1({ S6086, new_datapath_multdivunit_outmdu1_13 }),
  .out1({ S5143 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5557_ (
  .in1({ S6215, new_datapath_databusin_13 }),
  .out1({ S5144 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5558_ (
  .in1({ S5144, S5134 }),
  .out1({ S5145 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5559_ (
  .in1({ S5143, S5142 }),
  .out1({ S5146 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5560_ (
  .in1({ S5146, S5141 }),
  .out1({ S5148 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5561_ (
  .in1({ S5148, S5137 }),
  .out1({ S5149 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5562_ (
  .in1({ S5149, S5135 }),
  .out1({ S5150 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5563_ (
  .in1({ S5150, S5133 }),
  .out1({ S5151 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5564_ (
  .in1({ S5151, S5145 }),
  .out1({ S5152 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5565_ (
  .in1({ S5152, S5132 }),
  .out1({ S5153 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5566_ (
  .in1({ S5153, S5127 }),
  .out1({ S5154 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5567_ (
  .in1({ S5154, S5120 }),
  .out1({ new_datapath_indatatrf_13 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5568_ (
  .in1({ S5117, S4554 }),
  .out1({ S5155 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5569_ (
  .in1({ S5155, S4409 }),
  .out1({ S5156 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5570_ (
  .in1({ S5155, S4409 }),
  .out1({ S5158 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5571_ (
  .in1({ S5158, S4623 }),
  .out1({ S5159 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5572_ (
  .in1({ S5159, S5156 }),
  .out1({ S5160 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5573_ (
  .in1({ S5121, S4415 }),
  .out1({ S5161 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5574_ (
  .in1({ S5161, S4416 }),
  .out1({ S5162 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5575_ (
  .in1({ S5162, S4409 }),
  .out1({ S5163 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5576_ (
  .in1({ S5162, S4409 }),
  .out1({ S5164 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5577_ (
  .in1({ S5164, S4626 }),
  .out1({ S5165 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5578_ (
  .in1({ S5165, S5163 }),
  .out1({ S5166 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5579_ (
  .in1({ S5130, new_datapath_addsubunit_in1_14 }),
  .out1({ S5167 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5580_ (
  .in1({ S5129, S3390 }),
  .out1({ S5169 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5581_ (
  .in1({ S5169, S5167 }),
  .out1({ S5170 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5582_ (
  .in1({ S5170, S4637 }),
  .out1({ S5171 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5583_ (
  .in1({ S4660, new_datapath_shiftunit_2213_A }),
  .out1({ S5172 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5584_ (
  .in1({ S4648, new_datapath_shiftunit_2517_A }),
  .out1({ S5173 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5585_ (
  .in1({ S4629, S4408 }),
  .out1({ S5174 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5586_ (
  .in1({ S4285, new_controller_opcode_2 }),
  .out1({ S5175 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5587_ (
  .in1({ S5175, S4384 }),
  .out1({ S5176 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5588_ (
  .in1({ S5176, S4306 }),
  .out1({ S5177 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5589_ (
  .in1({ S5177, S4634 }),
  .out1({ S5178 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5590_ (
  .in1({ S6086, new_datapath_multdivunit_outmdu1_14 }),
  .out1({ S5180 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5591_ (
  .in1({ S3740, S3106 }),
  .out1({ S5181 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5592_ (
  .in1({ S4144, new_datapath_multdivunit_outmdu2_14 }),
  .out1({ S5182 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5593_ (
  .in1({ S5182, S5180 }),
  .out1({ S5183 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5594_ (
  .in1({ S5183, S5178 }),
  .out1({ S5184 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5595_ (
  .in1({ S5184, S5174 }),
  .out1({ S5185 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5596_ (
  .in1({ S5185, S5181 }),
  .out1({ S5186 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5597_ (
  .in1({ S5186, S5173 }),
  .out1({ S5187 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5598_ (
  .in1({ S4669, S161 }),
  .out1({ S5188 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5599_ (
  .in1({ S5188, S5172 }),
  .out1({ S5189 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5600_ (
  .in1({ S5189, S5187 }),
  .out1({ S5191 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5601_ (
  .in1({ S5191, S5171 }),
  .out1({ S5192 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5602_ (
  .in1({ S5192, S5160 }),
  .out1({ S5193 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5603_ (
  .in1({ S5193, S5166 }),
  .out1({ new_datapath_indatatrf_14 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5604_ (
  .in1({ S5158, S4406 }),
  .out1({ S5194 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5605_ (
  .in1({ S5194, S4401 }),
  .out1({ S5195 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5606_ (
  .in1({ S5194, S4401 }),
  .out1({ S5196 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5607_ (
  .in1({ S5196, S4624 }),
  .out1({ S5197 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5608_ (
  .in1({ S5197, S5195 }),
  .out1({ S5198 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5609_ (
  .in1({ S5164, S4408 }),
  .out1({ S5199 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5610_ (
  .in1({ S5199, S4401 }),
  .out1({ S5201 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5611_ (
  .in1({ S5199, S4401 }),
  .out1({ S5202 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5612_ (
  .in1({ S5201, S4625 }),
  .out1({ S5203 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5613_ (
  .in1({ S5203, S5202 }),
  .out1({ S5204 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5614_ (
  .in1({ S4670, S6075 }),
  .out1({ S5205 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5615_ (
  .in1({ S4660, new_datapath_shiftunit_2231_A }),
  .out1({ S5206 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5616_ (
  .in1({ S4648, new_datapath_shiftunit_2534_A }),
  .out1({ S5207 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5617_ (
  .in1({ S4629, new_datapath_addsubunit_in1_15 }),
  .out1({ S5208 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5618_ (
  .in1({ S5208, S4394 }),
  .out1({ S5209 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5619_ (
  .in1({ S4383, S4306 }),
  .out1({ S5210 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5620_ (
  .in1({ S5210, S4634 }),
  .out1({ S5212 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5621_ (
  .in1({ S4155, S2581 }),
  .out1({ S5213 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5622_ (
  .in1({ S3740, S2603 }),
  .out1({ S5214 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5623_ (
  .in1({ S6086, new_datapath_multdivunit_outmdu1_15 }),
  .out1({ S5215 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5624_ (
  .in1({ S5213, S5212 }),
  .out1({ S5216 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5625_ (
  .in1({ S5216, S5206 }),
  .out1({ S5217 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5626_ (
  .in1({ S5214, S5205 }),
  .out1({ S5218 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5627_ (
  .in1({ S5215, S5207 }),
  .out1({ S5219 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5628_ (
  .in1({ S5219, S5209 }),
  .out1({ S5220 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5629_ (
  .in1({ S5220, S5218 }),
  .out1({ S5221 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5630_ (
  .in1({ S5221, S5217 }),
  .out1({ S5223 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5631_ (
  .in1({ S5167, S3401 }),
  .out1({ S5224 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5632_ (
  .in1({ S5167, S3401 }),
  .out1({ S5225 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5633_ (
  .in1({ S5225, S4638 }),
  .out1({ S5226 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5634_ (
  .in1({ S5226, S5224 }),
  .out1({ S5227 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5635_ (
  .in1({ S5227, S5223 }),
  .out1({ S5228 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5636_ (
  .in1({ S5228, S5204 }),
  .out1({ S5229 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5637_ (
  .in1({ S5229, S5198 }),
  .out1({ new_datapath_indatatrf_15 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5638_ (
  .in1({ new_controller_1133_S_0, new_datapath_muxmem_in2_0 }),
  .out1({ S5230 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5639_ (
  .in1({ S3708, new_datapath_adr_outreg_0 }),
  .out1({ S5231 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5640_ (
  .in1({ S5231, S5230 }),
  .out1({ new_datapath_addrbus_0 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5641_ (
  .in1({ new_controller_1133_S_0, new_datapath_muxmem_in2_1 }),
  .out1({ S5233 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5642_ (
  .in1({ S3708, new_datapath_adr_outreg_1 }),
  .out1({ S5234 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5643_ (
  .in1({ S5234, S5233 }),
  .out1({ new_datapath_addrbus_1 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5644_ (
  .in1({ new_controller_1133_S_0, new_datapath_muxmem_in2_2 }),
  .out1({ S5235 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5645_ (
  .in1({ S3708, new_datapath_adr_outreg_2 }),
  .out1({ S5236 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5646_ (
  .in1({ S5236, S5235 }),
  .out1({ new_datapath_addrbus_2 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5647_ (
  .in1({ new_controller_1133_S_0, new_datapath_muxmem_in2_3 }),
  .out1({ S5237 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5648_ (
  .in1({ S3708, new_datapath_adr_outreg_3 }),
  .out1({ S5238 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5649_ (
  .in1({ S5238, S5237 }),
  .out1({ new_datapath_addrbus_3 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5650_ (
  .in1({ new_controller_1133_S_0, new_datapath_muxmem_in2_4 }),
  .out1({ S5240 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5651_ (
  .in1({ S3708, new_datapath_adr_outreg_4 }),
  .out1({ S5241 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5652_ (
  .in1({ S5241, S5240 }),
  .out1({ new_datapath_addrbus_4 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5653_ (
  .in1({ new_controller_1133_S_0, new_datapath_muxmem_in2_5 }),
  .out1({ S5242 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5654_ (
  .in1({ S3708, new_datapath_adr_outreg_5 }),
  .out1({ S5243 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5655_ (
  .in1({ S5243, S5242 }),
  .out1({ new_datapath_addrbus_5 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5656_ (
  .in1({ new_controller_1133_S_0, new_datapath_muxmem_in2_6 }),
  .out1({ S5244 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5657_ (
  .in1({ S3708, new_datapath_adr_outreg_6 }),
  .out1({ S5245 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5658_ (
  .in1({ S5245, S5244 }),
  .out1({ new_datapath_addrbus_6 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5659_ (
  .in1({ new_controller_1133_S_0, new_datapath_muxmem_in2_7 }),
  .out1({ S5246 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5660_ (
  .in1({ S3708, new_datapath_adr_outreg_7 }),
  .out1({ S5248 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5661_ (
  .in1({ S5248, S5246 }),
  .out1({ new_datapath_addrbus_7 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5662_ (
  .in1({ new_controller_1133_S_0, new_datapath_muxmem_in2_8 }),
  .out1({ S5249 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5663_ (
  .in1({ S3708, new_datapath_adr_outreg_8 }),
  .out1({ S5250 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5664_ (
  .in1({ S5250, S5249 }),
  .out1({ new_datapath_addrbus_8 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5665_ (
  .in1({ new_controller_1133_S_0, new_datapath_muxmem_in2_9 }),
  .out1({ S5251 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5666_ (
  .in1({ S3708, new_datapath_adr_outreg_9 }),
  .out1({ S5252 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5667_ (
  .in1({ S5252, S5251 }),
  .out1({ new_datapath_addrbus_9 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5668_ (
  .in1({ new_controller_1133_S_0, new_datapath_muxmem_in2_10 }),
  .out1({ S5253 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5669_ (
  .in1({ S3708, new_datapath_adr_outreg_10 }),
  .out1({ S5254 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5670_ (
  .in1({ S5254, S5253 }),
  .out1({ new_datapath_addrbus_10 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5671_ (
  .in1({ new_controller_1133_S_0, new_datapath_muxmem_in2_11 }),
  .out1({ S5256 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5672_ (
  .in1({ S3708, new_datapath_adr_outreg_11 }),
  .out1({ S5257 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5673_ (
  .in1({ S5257, S5256 }),
  .out1({ new_datapath_addrbus_11 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5674_ (
  .in1({ new_controller_1133_S_0, new_datapath_muxmem_in2_12 }),
  .out1({ S5258 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5675_ (
  .in1({ S3708, new_datapath_adr_outreg_12 }),
  .out1({ S5259 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5676_ (
  .in1({ S5259, S5258 }),
  .out1({ new_datapath_addrbus_12 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5677_ (
  .in1({ new_controller_1133_S_0, new_datapath_muxmem_in2_13 }),
  .out1({ S5260 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5678_ (
  .in1({ S3708, new_datapath_adr_outreg_13 }),
  .out1({ S5261 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5679_ (
  .in1({ S5261, S5260 }),
  .out1({ new_datapath_addrbus_13 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5680_ (
  .in1({ new_controller_1133_S_0, new_datapath_muxmem_in2_14 }),
  .out1({ S5263 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5681_ (
  .in1({ S3708, new_datapath_adr_outreg_14 }),
  .out1({ S5264 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5682_ (
  .in1({ S5264, S5263 }),
  .out1({ new_datapath_addrbus_14 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5683_ (
  .in1({ new_controller_1133_S_0, new_datapath_muxmem_in2_15 }),
  .out1({ S5265 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5684_ (
  .in1({ S3708, new_datapath_adr_outreg_15 }),
  .out1({ S5266 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5685_ (
  .in1({ S5266, S5265 }),
  .out1({ new_datapath_addrbus_15 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5686_ (
  .in1({ S6086, S6215 }),
  .out1({ S5267 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5687_ (
  .in1({ S5267, S4610 }),
  .out1({ S5268 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5688_ (
  .in1({ S5268 }),
  .out1({ S5269 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5689_ (
  .in1({ S5268, new_datapath_instruction_0 }),
  .out1({ S5270 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5690_ (
  .in1({ S4144, S2964 }),
  .out1({ S5272 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5691_ (
  .in1({ S5272, S5270 }),
  .out1({ new_datapath_muxrd_outmux_0 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5692_ (
  .in1({ new_datapath_instruction_1, new_datapath_instruction_0 }),
  .out1({ S5273 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5693_ (
  .in1({ S5268, new_datapath_instruction_1 }),
  .out1({ S5274 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5694_ (
  .in1({ new_datapath_instruction_1, new_datapath_instruction_0 }),
  .out1({ S5275 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5695_ (
  .in1({ S5275 }),
  .out1({ S5276 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5696_ (
  .in1({ S5273, S4155 }),
  .out1({ S5277 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5697_ (
  .in1({ S5277, S5275 }),
  .out1({ S5278 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5698_ (
  .in1({ S5278, S5274 }),
  .out1({ new_datapath_muxrd_outmux_1 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5699_ (
  .in1({ S5276, new_datapath_instruction_2 }),
  .out1({ S5279 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5700_ (
  .in1({ S5279, S4144 }),
  .out1({ S5281 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5701_ (
  .in1({ S5281 }),
  .out1({ S5282 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5702_ (
  .in1({ S5282, S5268 }),
  .out1({ S5283 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5703_ (
  .in1({ S5281, S5269 }),
  .out1({ S5284 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5704_ (
  .in1({ S5281, S5275 }),
  .out1({ S5285 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5705_ (
  .in1({ S5285, new_datapath_instruction_2 }),
  .out1({ S5286 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5706_ (
  .in1({ S5286, S5283 }),
  .out1({ new_datapath_muxrd_outmux_2 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5707_ (
  .in1({ S5279, S4155 }),
  .out1({ S5287 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5708_ (
  .in1({ S5287, new_datapath_instruction_3 }),
  .out1({ S5288 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5709_ (
  .in1({ S5284, S2975 }),
  .out1({ S5289 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5710_ (
  .in1({ S5289, S5288 }),
  .out1({ new_datapath_muxrd_outmux_3 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5711_ (
  .in1({ S270, S5693 }),
  .out1({ S5291 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5712_ (
  .in1({ S271, S5683 }),
  .out1({ S5292 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5713_ (
  .in1({ S5125, S2985 }),
  .out1({ S5293 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5714_ (
  .in1({ S5115, new_controller_fib_0 }),
  .out1({ S5294 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5715_ (
  .in1({ S5293, S5291 }),
  .out1({ S5295 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5716_ (
  .in1({ S5294, S5292 }),
  .out1({ S5296 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5717_ (
  .in1({ S256, S5693 }),
  .out1({ S5297 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5718_ (
  .in1({ S257, S5683 }),
  .out1({ S5298 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5719_ (
  .in1({ S5125, S3007 }),
  .out1({ S5299 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5720_ (
  .in1({ S5115, new_controller_fib_2 }),
  .out1({ S5301 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5721_ (
  .in1({ S5299, S5297 }),
  .out1({ S5302 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5722_ (
  .in1({ S5301, S5298 }),
  .out1({ S5303 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5723_ (
  .in1({ S264, S5693 }),
  .out1({ S5304 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5724_ (
  .in1({ S265, S5683 }),
  .out1({ S5305 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5725_ (
  .in1({ S5125, S2996 }),
  .out1({ S5306 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5726_ (
  .in1({ S5115, new_controller_fib_1 }),
  .out1({ S5307 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5727_ (
  .in1({ S5306, S5304 }),
  .out1({ S5308 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5728_ (
  .in1({ S5307, S5305 }),
  .out1({ S5309 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5729_ (
  .in1({ S248, S5693 }),
  .out1({ S5310 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5730_ (
  .in1({ S249, S5683 }),
  .out1({ S5312 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5731_ (
  .in1({ S5125, S3018 }),
  .out1({ S5313 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5732_ (
  .in1({ S5115, new_controller_fib_3 }),
  .out1({ S5314 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5733_ (
  .in1({ S5313, S5310 }),
  .out1({ S5315 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5734_ (
  .in1({ S5314, S5312 }),
  .out1({ S5316 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5735_ (
  .in1({ S5316, S5303 }),
  .out1({ S5317 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5736_ (
  .in1({ S5315, S5302 }),
  .out1({ S5318 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5737_ (
  .in1({ S5318, S5309 }),
  .out1({ S5319 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5738_ (
  .in1({ S5309, S5296 }),
  .out1({ S5320 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5739_ (
  .in1({ S5308, S5295 }),
  .out1({ S5321 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5740_ (
  .in1({ S5321, S5318 }),
  .out1({ S5323 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5741_ (
  .in1({ S5320, S5317 }),
  .out1({ S5324 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5742_ (
  .in1({ S5323, new_datapath_addsubunit_in1_0 }),
  .out1({ S5325 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5743_ (
  .in1({ S5325 }),
  .out1({ new_datapath_shiftunit_2265_A })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5744_ (
  .in1({ S5315, S5303 }),
  .out1({ S5326 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5745_ (
  .in1({ S5316, S5302 }),
  .out1({ S5327 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5746_ (
  .in1({ S5327, S5321 }),
  .out1({ S5328 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5747_ (
  .in1({ S5326, S5320 }),
  .out1({ S5329 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5748_ (
  .in1({ S5328, new_datapath_addsubunit_in1_8 }),
  .out1({ S5330 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5749_ (
  .in1({ S5308, S5295 }),
  .out1({ S5331 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5750_ (
  .in1({ S5309, S5296 }),
  .out1({ S5333 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5751_ (
  .in1({ S5316, S5302 }),
  .out1({ S5334 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5752_ (
  .in1({ S5315, S5303 }),
  .out1({ S5335 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5753_ (
  .in1({ S5335, S5333 }),
  .out1({ S5336 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5754_ (
  .in1({ S5334, S5331 }),
  .out1({ S5337 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5755_ (
  .in1({ S5336, new_datapath_addsubunit_in1_7 }),
  .out1({ S5338 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5756_ (
  .in1({ S5309, S5295 }),
  .out1({ S5339 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5757_ (
  .in1({ S5308, S5296 }),
  .out1({ S5340 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5758_ (
  .in1({ S5315, S5302 }),
  .out1({ S5341 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5759_ (
  .in1({ S5316, S5303 }),
  .out1({ S5342 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5760_ (
  .in1({ S5342, S5340 }),
  .out1({ S5344 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5761_ (
  .in1({ S5344, new_datapath_addsubunit_in1_13 }),
  .out1({ S5345 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5762_ (
  .in1({ S5340, S5327 }),
  .out1({ S5346 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5763_ (
  .in1({ S5346, new_datapath_addsubunit_in1_9 }),
  .out1({ S5347 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5764_ (
  .in1({ S5347, S5345 }),
  .out1({ S5348 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5765_ (
  .in1({ S5340, S5335 }),
  .out1({ S5349 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5766_ (
  .in1({ S5349, new_datapath_addsubunit_in1_5 }),
  .out1({ S5350 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5767_ (
  .in1({ S5342, S3401 }),
  .out1({ S5351 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5768_ (
  .in1({ S5351, S5331 }),
  .out1({ S5352 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5769_ (
  .in1({ S5333, S5327 }),
  .out1({ S5353 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5770_ (
  .in1({ S5353, new_datapath_addsubunit_in1_11 }),
  .out1({ S5355 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5771_ (
  .in1({ S5308, S5296 }),
  .out1({ S5356 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5772_ (
  .in1({ S5309, S5295 }),
  .out1({ S5357 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5773_ (
  .in1({ S5357, S5342 }),
  .out1({ S5358 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5774_ (
  .in1({ S5358, new_datapath_addsubunit_in1_14 }),
  .out1({ S5359 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5775_ (
  .in1({ S5342, S5321 }),
  .out1({ S5360 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5776_ (
  .in1({ S5341, S5320 }),
  .out1({ S5361 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5777_ (
  .in1({ S5360, new_datapath_addsubunit_in1_12 }),
  .out1({ S5362 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5778_ (
  .in1({ S5335, S5321 }),
  .out1({ S5363 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5779_ (
  .in1({ S5334, S5320 }),
  .out1({ S5364 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5780_ (
  .in1({ S5363, new_datapath_addsubunit_in1_4 }),
  .out1({ S5366 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5781_ (
  .in1({ S5333, S5318 }),
  .out1({ S5367 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5782_ (
  .in1({ S5331, S5317 }),
  .out1({ S5368 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5783_ (
  .in1({ S5367, new_datapath_addsubunit_in1_3 }),
  .out1({ S5369 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5784_ (
  .in1({ S5357, S5335 }),
  .out1({ S5370 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5785_ (
  .in1({ S5370, new_datapath_addsubunit_in1_6 }),
  .out1({ S5371 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5786_ (
  .in1({ S5357, S5318 }),
  .out1({ S5372 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5787_ (
  .in1({ S5356, S5317 }),
  .out1({ S5373 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5788_ (
  .in1({ S5372, new_datapath_addsubunit_in1_2 }),
  .out1({ S5374 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5789_ (
  .in1({ S5357, S5327 }),
  .out1({ S5375 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5790_ (
  .in1({ S5375, new_datapath_addsubunit_in1_10 }),
  .out1({ S5377 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5791_ (
  .in1({ S5369, S5325 }),
  .out1({ S5378 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5792_ (
  .in1({ S5371, S5350 }),
  .out1({ S5379 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5793_ (
  .in1({ S5379, S5378 }),
  .out1({ S5380 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5794_ (
  .in1({ S5377, S5355 }),
  .out1({ S5381 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5795_ (
  .in1({ S5362, S5359 }),
  .out1({ S5382 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5796_ (
  .in1({ S5382, S5381 }),
  .out1({ S5383 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5797_ (
  .in1({ S5383, S5380 }),
  .out1({ S5384 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5798_ (
  .in1({ S5366, S5330 }),
  .out1({ S5385 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5799_ (
  .in1({ S5385, S5348 }),
  .out1({ S5386 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5800_ (
  .in1({ S5374, S5352 }),
  .out1({ S5388 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5801_ (
  .in1({ S5340, S5318 }),
  .out1({ S5389 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5802_ (
  .in1({ S5339, S5317 }),
  .out1({ S5390 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5803_ (
  .in1({ S5390, S5966 }),
  .out1({ S5391 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5804_ (
  .in1({ S5389, new_datapath_addsubunit_in1_1 }),
  .out1({ S5392 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5805_ (
  .in1({ S5392, S5338 }),
  .out1({ S5393 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5806_ (
  .in1({ S5393, S5388 }),
  .out1({ S5394 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5807_ (
  .in1({ S5394, S5386 }),
  .out1({ S5395 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5808_ (
  .in1({ S5342, S5333 }),
  .out1({ S5396 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5809_ (
  .in1({ S5395, S5384 }),
  .out1({ S5397 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5810_ (
  .in1({ S5397 }),
  .out1({ new_datapath_shiftunit_1961_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5811_ (
  .in1({ S5323, new_datapath_addsubunit_in1_1 }),
  .out1({ S5399 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5812_ (
  .in1({ S5363, new_datapath_addsubunit_in1_5 }),
  .out1({ S5400 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5813_ (
  .in1({ S5360, new_datapath_addsubunit_in1_13 }),
  .out1({ S5401 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5814_ (
  .in1({ S5356, S5351 }),
  .out1({ S5402 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5815_ (
  .in1({ S5353, new_datapath_addsubunit_in1_12 }),
  .out1({ S5403 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5816_ (
  .in1({ S5370, new_datapath_addsubunit_in1_7 }),
  .out1({ S5404 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5817_ (
  .in1({ S5349, new_datapath_addsubunit_in1_6 }),
  .out1({ S5405 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5818_ (
  .in1({ S5336, new_datapath_addsubunit_in1_8 }),
  .out1({ S5406 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5819_ (
  .in1({ S5406 }),
  .out1({ S5407 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5820_ (
  .in1({ S5375, new_datapath_addsubunit_in1_11 }),
  .out1({ S5409 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5821_ (
  .in1({ S5372, new_datapath_addsubunit_in1_3 }),
  .out1({ S5410 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5822_ (
  .in1({ S5367, new_datapath_addsubunit_in1_4 }),
  .out1({ S5411 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5823_ (
  .in1({ S5344, new_datapath_addsubunit_in1_14 }),
  .out1({ S5412 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5824_ (
  .in1({ S5412 }),
  .out1({ S5413 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5825_ (
  .in1({ S5346, new_datapath_addsubunit_in1_10 }),
  .out1({ S5414 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5826_ (
  .in1({ S5328, new_datapath_addsubunit_in1_9 }),
  .out1({ S5415 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5827_ (
  .in1({ S5414, S5410 }),
  .out1({ S5416 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5828_ (
  .in1({ S5401, S5399 }),
  .out1({ S5417 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5829_ (
  .in1({ S5417, S5416 }),
  .out1({ S5418 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5830_ (
  .in1({ S5390, S5957 }),
  .out1({ S5420 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5831_ (
  .in1({ S4652, S3401 }),
  .out1({ S5421 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5832_ (
  .in1({ S4653, new_datapath_addsubunit_in1_15 }),
  .out1({ S5422 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5833_ (
  .in1({ S5422, S5315 }),
  .out1({ S5423 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5834_ (
  .in1({ S5421, S5341 }),
  .out1({ S5424 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5835_ (
  .in1({ S5424 }),
  .out1({ S5425 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5836_ (
  .in1({ S5424, S5333 }),
  .out1({ S5426 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5837_ (
  .in1({ S5426, S5420 }),
  .out1({ S5427 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5838_ (
  .in1({ S5409, S5400 }),
  .out1({ S5428 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5839_ (
  .in1({ S5428, S5407 }),
  .out1({ S5429 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5840_ (
  .in1({ S5429, S5427 }),
  .out1({ S5431 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5841_ (
  .in1({ S5415, S5402 }),
  .out1({ S5432 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5842_ (
  .in1({ S5432, S5413 }),
  .out1({ S5433 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5843_ (
  .in1({ S5411, S5404 }),
  .out1({ S5434 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5844_ (
  .in1({ S5405, S5403 }),
  .out1({ S5435 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5845_ (
  .in1({ S5435, S5434 }),
  .out1({ S5436 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5846_ (
  .in1({ S5436, S5433 }),
  .out1({ S5437 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5847_ (
  .in1({ S5437, S5431 }),
  .out1({ S5438 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5848_ (
  .in1({ S5438, S5418 }),
  .out1({ new_datapath_shiftunit_1979_A })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5849_ (
  .in1({ S5324, S5957 }),
  .out1({ S5439 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5850_ (
  .in1({ S5323, new_datapath_addsubunit_in1_2 }),
  .out1({ S5441 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5851_ (
  .in1({ S5372, new_datapath_addsubunit_in1_4 }),
  .out1({ S5442 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5852_ (
  .in1({ S5328, new_datapath_addsubunit_in1_10 }),
  .out1({ S5443 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5853_ (
  .in1({ S5375, new_datapath_addsubunit_in1_12 }),
  .out1({ S5444 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5854_ (
  .in1({ S5349, new_datapath_addsubunit_in1_7 }),
  .out1({ S5445 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5855_ (
  .in1({ S5370, new_datapath_addsubunit_in1_8 }),
  .out1({ S5446 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5856_ (
  .in1({ S5360, new_datapath_addsubunit_in1_14 }),
  .out1({ S5447 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5857_ (
  .in1({ S5353, new_datapath_addsubunit_in1_13 }),
  .out1({ S5448 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5858_ (
  .in1({ S5346, new_datapath_addsubunit_in1_11 }),
  .out1({ S5449 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5859_ (
  .in1({ S5336, new_datapath_addsubunit_in1_9 }),
  .out1({ S5450 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5860_ (
  .in1({ S5423, S5309 }),
  .out1({ S5452 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5861_ (
  .in1({ S5367, new_datapath_addsubunit_in1_5 }),
  .out1({ S5453 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5862_ (
  .in1({ S5364, S5916 }),
  .out1({ S5454 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5863_ (
  .in1({ S5363, new_datapath_addsubunit_in1_6 }),
  .out1({ S5455 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5864_ (
  .in1({ S5344, new_datapath_addsubunit_in1_15 }),
  .out1({ S5456 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5865_ (
  .in1({ S5456, S5450 }),
  .out1({ S5457 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5866_ (
  .in1({ S5457, S5439 }),
  .out1({ S5458 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5867_ (
  .in1({ S5453, S5445 }),
  .out1({ S5459 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5868_ (
  .in1({ S5425, S5309 }),
  .out1({ S5460 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5869_ (
  .in1({ S5460, S5447 }),
  .out1({ S5461 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5870_ (
  .in1({ S5461, S5459 }),
  .out1({ S5463 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5871_ (
  .in1({ S5463, S5458 }),
  .out1({ S5464 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5872_ (
  .in1({ S5448, S5443 }),
  .out1({ S5465 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5873_ (
  .in1({ S5389, new_datapath_addsubunit_in1_3 }),
  .out1({ S5466 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5874_ (
  .in1({ S5466, S5444 }),
  .out1({ S5467 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5875_ (
  .in1({ S5467, S5465 }),
  .out1({ S5468 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5876_ (
  .in1({ S5449, S5442 }),
  .out1({ S5469 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5877_ (
  .in1({ S5455, S5446 }),
  .out1({ S5470 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5878_ (
  .in1({ S5470, S5469 }),
  .out1({ S5471 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5879_ (
  .in1({ S5471, S5468 }),
  .out1({ S5472 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5880_ (
  .in1({ S5472, S5464 }),
  .out1({ S5474 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5881_ (
  .in1({ S5474 }),
  .out1({ new_datapath_shiftunit_1997_A })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5882_ (
  .in1({ S5364, S5907 }),
  .out1({ S5475 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5883_ (
  .in1({ S5363, new_datapath_addsubunit_in1_7 }),
  .out1({ S5476 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5884_ (
  .in1({ S5367, new_datapath_addsubunit_in1_6 }),
  .out1({ S5477 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5885_ (
  .in1({ S5353, new_datapath_addsubunit_in1_14 }),
  .out1({ S5478 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5886_ (
  .in1({ S5336, new_datapath_addsubunit_in1_10 }),
  .out1({ S5479 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5887_ (
  .in1({ S5479 }),
  .out1({ S5480 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5888_ (
  .in1({ S5324, S5947 }),
  .out1({ S5481 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5889_ (
  .in1({ S5328, new_datapath_addsubunit_in1_11 }),
  .out1({ S5482 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5890_ (
  .in1({ S5482 }),
  .out1({ S5484 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5891_ (
  .in1({ S5346, new_datapath_addsubunit_in1_12 }),
  .out1({ S5485 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5892_ (
  .in1({ S5370, new_datapath_addsubunit_in1_9 }),
  .out1({ S5486 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5893_ (
  .in1({ S5321, S4652 }),
  .out1({ S5487 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5894_ (
  .in1({ S5487, S5351 }),
  .out1({ S5488 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5895_ (
  .in1({ S5349, new_datapath_addsubunit_in1_8 }),
  .out1({ S5489 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5896_ (
  .in1({ S5372, new_datapath_addsubunit_in1_5 }),
  .out1({ S5490 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5897_ (
  .in1({ S5375, new_datapath_addsubunit_in1_13 }),
  .out1({ S5491 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5898_ (
  .in1({ S5491, S5485 }),
  .out1({ S5492 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5899_ (
  .in1({ S5492, S5484 }),
  .out1({ S5493 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5900_ (
  .in1({ S5493, S5488 }),
  .out1({ S5495 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5901_ (
  .in1({ S5490, S5478 }),
  .out1({ S5496 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5902_ (
  .in1({ S5389, new_datapath_addsubunit_in1_4 }),
  .out1({ S5497 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5903_ (
  .in1({ S5496, S5475 }),
  .out1({ S5498 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5904_ (
  .in1({ S5481, S5480 }),
  .out1({ S5499 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5905_ (
  .in1({ S5497, S5477 }),
  .out1({ S5500 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5906_ (
  .in1({ S5489, S5486 }),
  .out1({ S5501 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5907_ (
  .in1({ S5501, S5500 }),
  .out1({ S5502 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5908_ (
  .in1({ S5502, S5499 }),
  .out1({ S5503 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5909_ (
  .in1({ S5503, S5495 }),
  .out1({ S5504 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5910_ (
  .in1({ S5504, S5498 }),
  .out1({ new_datapath_shiftunit_2015_A })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5911_ (
  .in1({ S5324, S5936 }),
  .out1({ S5506 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5912_ (
  .in1({ S5323, new_datapath_addsubunit_in1_4 }),
  .out1({ S5507 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5913_ (
  .in1({ S5390, S5926 }),
  .out1({ S5508 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5914_ (
  .in1({ S5389, new_datapath_addsubunit_in1_5 }),
  .out1({ S5509 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5915_ (
  .in1({ S5508, S5506 }),
  .out1({ S5510 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5916_ (
  .in1({ S5375, new_datapath_addsubunit_in1_14 }),
  .out1({ S5511 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5917_ (
  .in1({ S5363, new_datapath_addsubunit_in1_8 }),
  .out1({ S5512 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5918_ (
  .in1({ S5349, new_datapath_addsubunit_in1_9 }),
  .out1({ S5513 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5919_ (
  .in1({ S5513 }),
  .out1({ S5514 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5920_ (
  .in1({ S5370, new_datapath_addsubunit_in1_10 }),
  .out1({ S5516 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5921_ (
  .in1({ S5373, S5916 }),
  .out1({ S5517 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5922_ (
  .in1({ S5328, new_datapath_addsubunit_in1_12 }),
  .out1({ S5518 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5923_ (
  .in1({ S5353, new_datapath_addsubunit_in1_15 }),
  .out1({ S5519 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5924_ (
  .in1({ S5368, S5907 }),
  .out1({ S5520 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5925_ (
  .in1({ S5367, new_datapath_addsubunit_in1_7 }),
  .out1({ S5521 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5926_ (
  .in1({ S5336, new_datapath_addsubunit_in1_11 }),
  .out1({ S5522 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5927_ (
  .in1({ S5346, new_datapath_addsubunit_in1_13 }),
  .out1({ S5523 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5928_ (
  .in1({ S5520, S5517 }),
  .out1({ S5524 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5929_ (
  .in1({ S5522, S5511 }),
  .out1({ S5525 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5930_ (
  .in1({ S5523, S5512 }),
  .out1({ S5527 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5931_ (
  .in1({ S5519, S5424 }),
  .out1({ S5528 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5932_ (
  .in1({ S5528, S5527 }),
  .out1({ S5529 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5933_ (
  .in1({ S5529 }),
  .out1({ S5530 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5934_ (
  .in1({ S5530, S5525 }),
  .out1({ S5531 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5935_ (
  .in1({ S5524, S5510 }),
  .out1({ S5532 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5936_ (
  .in1({ S5518, S5513 }),
  .out1({ S5533 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5937_ (
  .in1({ S5533 }),
  .out1({ S5534 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5938_ (
  .in1({ S5534, S5516 }),
  .out1({ S5535 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5939_ (
  .in1({ S5535, S5532 }),
  .out1({ S5536 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5940_ (
  .in1({ S5536, S5531 }),
  .out1({ new_datapath_shiftunit_2033_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5941_ (
  .in1({ S5367, new_datapath_addsubunit_in1_8 }),
  .out1({ S5538 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5942_ (
  .in1({ S5349, new_datapath_addsubunit_in1_10 }),
  .out1({ S5539 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5943_ (
  .in1({ S5421, S5353 }),
  .out1({ S5540 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5944_ (
  .in1({ S5323, new_datapath_addsubunit_in1_5 }),
  .out1({ S5541 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5945_ (
  .in1({ S5363, new_datapath_addsubunit_in1_9 }),
  .out1({ S5542 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5946_ (
  .in1({ S5372, new_datapath_addsubunit_in1_7 }),
  .out1({ S5543 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5947_ (
  .in1({ S5328, new_datapath_addsubunit_in1_13 }),
  .out1({ S5544 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5948_ (
  .in1({ S5544, S5543 }),
  .out1({ S5545 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5949_ (
  .in1({ S5370, new_datapath_addsubunit_in1_11 }),
  .out1({ S5546 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5950_ (
  .in1({ S5375, new_datapath_addsubunit_in1_15 }),
  .out1({ S5548 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5951_ (
  .in1({ S5336, new_datapath_addsubunit_in1_12 }),
  .out1({ S5549 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5952_ (
  .in1({ S5346, new_datapath_addsubunit_in1_14 }),
  .out1({ S5550 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5953_ (
  .in1({ S5546, S5542 }),
  .out1({ S5551 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5954_ (
  .in1({ S5551 }),
  .out1({ S5552 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5955_ (
  .in1({ S5552, S5549 }),
  .out1({ S5553 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5956_ (
  .in1({ S5548, S5538 }),
  .out1({ S5554 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5957_ (
  .in1({ S5554, S5545 }),
  .out1({ S5555 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5958_ (
  .in1({ S5555 }),
  .out1({ S5556 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5959_ (
  .in1({ S5556, S5553 }),
  .out1({ S5557 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5960_ (
  .in1({ S5539, S5424 }),
  .out1({ S5559 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5961_ (
  .in1({ S5389, new_datapath_addsubunit_in1_6 }),
  .out1({ S5560 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5962_ (
  .in1({ S5560, S5550 }),
  .out1({ S5561 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5963_ (
  .in1({ S5541, S5540 }),
  .out1({ S5562 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5964_ (
  .in1({ S5562, S5561 }),
  .out1({ S5563 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5965_ (
  .in1({ S5563 }),
  .out1({ S5564 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5966_ (
  .in1({ S5564, S5559 }),
  .out1({ S5565 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5967_ (
  .in1({ S5565, S5557 }),
  .out1({ new_datapath_shiftunit_2051_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5968_ (
  .in1({ S5336, new_datapath_addsubunit_in1_13 }),
  .out1({ S5566 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5969_ (
  .in1({ S5349, new_datapath_addsubunit_in1_11 }),
  .out1({ S5567 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5970_ (
  .in1({ S5567, S5566 }),
  .out1({ S5569 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5971_ (
  .in1({ S5323, new_datapath_addsubunit_in1_6 }),
  .out1({ S5570 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5972_ (
  .in1({ S5370, new_datapath_addsubunit_in1_12 }),
  .out1({ S5571 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5973_ (
  .in1({ S5363, new_datapath_addsubunit_in1_10 }),
  .out1({ S5572 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5974_ (
  .in1({ S5452, S5424 }),
  .out1({ S5573 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5975_ (
  .in1({ S5372, new_datapath_addsubunit_in1_8 }),
  .out1({ S5574 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5976_ (
  .in1({ S5328, new_datapath_addsubunit_in1_14 }),
  .out1({ S5575 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5977_ (
  .in1({ S5575, S5574 }),
  .out1({ S5576 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5978_ (
  .in1({ S5367, new_datapath_addsubunit_in1_9 }),
  .out1({ S5577 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5979_ (
  .in1({ S5346, new_datapath_addsubunit_in1_15 }),
  .out1({ S5578 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5980_ (
  .in1({ S5390, S5907 }),
  .out1({ S5580 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5981_ (
  .in1({ S5389, new_datapath_addsubunit_in1_7 }),
  .out1({ S5581 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5982_ (
  .in1({ S5581, S5571 }),
  .out1({ S5582 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5983_ (
  .in1({ S5582, S5569 }),
  .out1({ S5583 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5984_ (
  .in1({ S5578, S5570 }),
  .out1({ S5584 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5985_ (
  .in1({ S5577, S5572 }),
  .out1({ S5585 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5986_ (
  .in1({ S5585, S5584 }),
  .out1({ S5586 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_5987_ (
  .in1({ S5576, S5573 }),
  .out1({ S5587 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5988_ (
  .in1({ S5587, S5586 }),
  .out1({ S5588 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_5989_ (
  .in1({ S5588 }),
  .out1({ S5589 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5990_ (
  .in1({ S5589, S5583 }),
  .out1({ new_datapath_shiftunit_2069_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5991_ (
  .in1({ S5323, new_datapath_addsubunit_in1_7 }),
  .out1({ S5591 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5992_ (
  .in1({ S5421, S5346 }),
  .out1({ S5592 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5993_ (
  .in1({ S5328, new_datapath_addsubunit_in1_15 }),
  .out1({ S5593 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5994_ (
  .in1({ S5370, new_datapath_addsubunit_in1_13 }),
  .out1({ S5594 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5995_ (
  .in1({ S5372, new_datapath_addsubunit_in1_9 }),
  .out1({ S5595 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5996_ (
  .in1({ S5363, new_datapath_addsubunit_in1_11 }),
  .out1({ S5596 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5997_ (
  .in1({ S5349, new_datapath_addsubunit_in1_12 }),
  .out1({ S5597 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5998_ (
  .in1({ S5336, new_datapath_addsubunit_in1_14 }),
  .out1({ S5598 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_5999_ (
  .in1({ S5367, new_datapath_addsubunit_in1_10 }),
  .out1({ S5599 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6000_ (
  .in1({ S5389, new_datapath_addsubunit_in1_8 }),
  .out1({ S5601 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6001_ (
  .in1({ S5601, S5594 }),
  .out1({ S5602 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6002_ (
  .in1({ S5597, S5593 }),
  .out1({ S5603 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6003_ (
  .in1({ S5603, S5602 }),
  .out1({ S5604 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6004_ (
  .in1({ S5595, S5592 }),
  .out1({ S5605 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6005_ (
  .in1({ S5599, S5591 }),
  .out1({ S5606 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6006_ (
  .in1({ S5606, S5605 }),
  .out1({ S5607 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6007_ (
  .in1({ S5598, S5596 }),
  .out1({ S5608 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6008_ (
  .in1({ S5608, S5573 }),
  .out1({ S5609 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6009_ (
  .in1({ S5609, S5607 }),
  .out1({ S5610 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6010_ (
  .in1({ S5610 }),
  .out1({ S5612 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6011_ (
  .in1({ S5612, S5604 }),
  .out1({ new_datapath_shiftunit_2087_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6012_ (
  .in1({ S5349, new_datapath_addsubunit_in1_13 }),
  .out1({ S5613 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6013_ (
  .in1({ S5370, new_datapath_addsubunit_in1_14 }),
  .out1({ S5614 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6014_ (
  .in1({ S5336, new_datapath_addsubunit_in1_15 }),
  .out1({ S5615 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6015_ (
  .in1({ S5323, new_datapath_addsubunit_in1_8 }),
  .out1({ S5616 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6016_ (
  .in1({ S5389, new_datapath_addsubunit_in1_9 }),
  .out1({ S5617 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6017_ (
  .in1({ S5617, S5616 }),
  .out1({ S5618 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6018_ (
  .in1({ S5618 }),
  .out1({ S5619 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6019_ (
  .in1({ S5368, S3357 }),
  .out1({ S5620 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6020_ (
  .in1({ S5367, new_datapath_addsubunit_in1_11 }),
  .out1({ S5622 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6021_ (
  .in1({ S5620, S5423 }),
  .out1({ S5623 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6022_ (
  .in1({ S5363, new_datapath_addsubunit_in1_12 }),
  .out1({ S5624 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6023_ (
  .in1({ S5372, new_datapath_addsubunit_in1_10 }),
  .out1({ S5625 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6024_ (
  .in1({ S5625, S5624 }),
  .out1({ S5626 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6025_ (
  .in1({ S5614, S5613 }),
  .out1({ S5627 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6026_ (
  .in1({ S5627, S5626 }),
  .out1({ S5628 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6027_ (
  .in1({ S5628 }),
  .out1({ S5629 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6028_ (
  .in1({ S5619, S5615 }),
  .out1({ S5630 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6029_ (
  .in1({ S5630, S5629 }),
  .out1({ S5631 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6030_ (
  .in1({ S5631, S5623 }),
  .out1({ new_datapath_shiftunit_2105_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6031_ (
  .in1({ S5363, new_datapath_addsubunit_in1_13 }),
  .out1({ S5633 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6032_ (
  .in1({ S5372, new_datapath_addsubunit_in1_11 }),
  .out1({ S5634 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6033_ (
  .in1({ S5367, new_datapath_addsubunit_in1_12 }),
  .out1({ S5635 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6034_ (
  .in1({ S5349, new_datapath_addsubunit_in1_14 }),
  .out1({ S5636 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6035_ (
  .in1({ S5370, S4653 }),
  .out1({ S5637 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6036_ (
  .in1({ S5309, S5303 }),
  .out1({ S5638 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6037_ (
  .in1({ S5638 }),
  .out1({ S5639 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6038_ (
  .in1({ S5639, S5316 }),
  .out1({ S5640 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6039_ (
  .in1({ S5638, S5315 }),
  .out1({ S5641 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6040_ (
  .in1({ S5637, S3401 }),
  .out1({ S5643 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6041_ (
  .in1({ S5643, S5641 }),
  .out1({ S5644 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6042_ (
  .in1({ S5323, new_datapath_addsubunit_in1_9 }),
  .out1({ S5645 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6043_ (
  .in1({ S5645, S5644 }),
  .out1({ S5646 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6044_ (
  .in1({ S5389, new_datapath_addsubunit_in1_10 }),
  .out1({ S5647 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6045_ (
  .in1({ S5635, S5633 }),
  .out1({ S5648 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6046_ (
  .in1({ S5636, S5634 }),
  .out1({ S5649 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6047_ (
  .in1({ S5649, S5648 }),
  .out1({ S5650 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6048_ (
  .in1({ S5650, S5647 }),
  .out1({ S5651 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6049_ (
  .in1({ S5651, S5646 }),
  .out1({ S5652 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6050_ (
  .in1({ S5652 }),
  .out1({ new_datapath_shiftunit_2123_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6051_ (
  .in1({ S5349, new_datapath_addsubunit_in1_15 }),
  .out1({ S5654 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6052_ (
  .in1({ S5363, new_datapath_addsubunit_in1_14 }),
  .out1({ S5655 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6053_ (
  .in1({ S5655, S5654 }),
  .out1({ S5656 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6054_ (
  .in1({ S5372, new_datapath_addsubunit_in1_12 }),
  .out1({ S5657 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6055_ (
  .in1({ S5367, new_datapath_addsubunit_in1_13 }),
  .out1({ S5658 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6056_ (
  .in1({ S5323, new_datapath_addsubunit_in1_10 }),
  .out1({ S5659 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6057_ (
  .in1({ S5640, S5422 }),
  .out1({ S5660 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6058_ (
  .in1({ S5660, S5656 }),
  .out1({ S5661 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6059_ (
  .in1({ S5389, new_datapath_addsubunit_in1_11 }),
  .out1({ S5662 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6060_ (
  .in1({ S5662, S5657 }),
  .out1({ S5664 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6061_ (
  .in1({ S5659, S5658 }),
  .out1({ S5665 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6062_ (
  .in1({ S5665, S5664 }),
  .out1({ S5666 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6063_ (
  .in1({ S5666, S5661 }),
  .out1({ new_datapath_shiftunit_2141_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6064_ (
  .in1({ S5421, S5349 }),
  .out1({ S5667 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6065_ (
  .in1({ S5367, new_datapath_addsubunit_in1_14 }),
  .out1({ S5668 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6066_ (
  .in1({ S5668, S5667 }),
  .out1({ S5669 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6067_ (
  .in1({ S5372, new_datapath_addsubunit_in1_13 }),
  .out1({ S5670 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6068_ (
  .in1({ S5363, new_datapath_addsubunit_in1_15 }),
  .out1({ S5671 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6069_ (
  .in1({ S5323, new_datapath_addsubunit_in1_11 }),
  .out1({ S5672 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6070_ (
  .in1({ S5672, S5670 }),
  .out1({ S5674 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6071_ (
  .in1({ S5389, new_datapath_addsubunit_in1_12 }),
  .out1({ S5675 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6072_ (
  .in1({ S5675, S5671 }),
  .out1({ S5676 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6073_ (
  .in1({ S5676, S5674 }),
  .out1({ S5677 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6074_ (
  .in1({ S5669, S5660 }),
  .out1({ S5678 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6075_ (
  .in1({ S5678, S5677 }),
  .out1({ new_datapath_shiftunit_2159_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6076_ (
  .in1({ S5323, new_datapath_addsubunit_in1_12 }),
  .out1({ S5679 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6077_ (
  .in1({ S5372, new_datapath_addsubunit_in1_14 }),
  .out1({ S5680 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6078_ (
  .in1({ S5331, S5318 }),
  .out1({ S5681 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6079_ (
  .in1({ S5318, S4652 }),
  .out1({ S5682 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6080_ (
  .in1({ S5682, new_datapath_addsubunit_in1_15 }),
  .out1({ S5684 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6081_ (
  .in1({ S5684, S5681 }),
  .out1({ S5685 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6082_ (
  .in1({ S5389, new_datapath_addsubunit_in1_13 }),
  .out1({ S5686 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6083_ (
  .in1({ S5686, S5680 }),
  .out1({ S5687 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6084_ (
  .in1({ S5687, S5685 }),
  .out1({ S5688 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6085_ (
  .in1({ S5688, S5679 }),
  .out1({ new_datapath_shiftunit_2177_A })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6086_ (
  .in1({ S5681, S4652 }),
  .out1({ S5689 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6087_ (
  .in1({ S5689, S5372 }),
  .out1({ S5690 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6088_ (
  .in1({ S5690, S3401 }),
  .out1({ S5691 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6089_ (
  .in1({ S5323, new_datapath_addsubunit_in1_13 }),
  .out1({ S5692 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6090_ (
  .in1({ S5389, new_datapath_addsubunit_in1_14 }),
  .out1({ S5694 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6091_ (
  .in1({ S5694, S5692 }),
  .out1({ S5695 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6092_ (
  .in1({ S5695, S5691 }),
  .out1({ S5696 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6093_ (
  .in1({ S5696 }),
  .out1({ new_datapath_shiftunit_2195_A })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6094_ (
  .in1({ S5422, S5319 }),
  .out1({ S5697 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6095_ (
  .in1({ S5323, new_datapath_addsubunit_in1_14 }),
  .out1({ S5698 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6096_ (
  .in1({ S5389, new_datapath_addsubunit_in1_15 }),
  .out1({ S5699 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6097_ (
  .in1({ S5699 }),
  .out1({ S5700 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6098_ (
  .in1({ S5700, S5697 }),
  .out1({ S5701 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6099_ (
  .in1({ S5701, S5698 }),
  .out1({ new_datapath_shiftunit_2213_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6100_ (
  .in1({ S5323, new_datapath_addsubunit_in1_15 }),
  .out1({ S5703 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6101_ (
  .in1({ S5703, S5422 }),
  .out1({ new_datapath_shiftunit_2231_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6102_ (
  .in1({ S5389, new_datapath_addsubunit_in1_0 }),
  .out1({ S5704 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6103_ (
  .in1({ S5704, S5399 }),
  .out1({ new_datapath_shiftunit_2283_A })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6104_ (
  .in1({ S5373, S5975 }),
  .out1({ S5705 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6105_ (
  .in1({ S5705, S5391 }),
  .out1({ S5706 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6106_ (
  .in1({ S5706, S5441 }),
  .out1({ new_datapath_shiftunit_2301_A })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6107_ (
  .in1({ S5373, S5966 }),
  .out1({ S5707 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6108_ (
  .in1({ S5368, S5975 }),
  .out1({ S5708 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6109_ (
  .in1({ S5707, S5420 }),
  .out1({ S5709 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6110_ (
  .in1({ S5708, S5481 }),
  .out1({ S5711 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6111_ (
  .in1({ S5711, S5709 }),
  .out1({ new_datapath_shiftunit_2319_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6112_ (
  .in1({ S5367, new_datapath_addsubunit_in1_1 }),
  .out1({ S5712 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6113_ (
  .in1({ S5363, new_datapath_addsubunit_in1_0 }),
  .out1({ S5713 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6114_ (
  .in1({ S5712, S5507 }),
  .out1({ S5714 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6115_ (
  .in1({ S5466, S5374 }),
  .out1({ S5715 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6116_ (
  .in1({ S5715, S5714 }),
  .out1({ S5716 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6117_ (
  .in1({ S5716, S5713 }),
  .out1({ new_datapath_shiftunit_2337_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6118_ (
  .in1({ S5367, new_datapath_addsubunit_in1_2 }),
  .out1({ S5717 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6119_ (
  .in1({ S5349, new_datapath_addsubunit_in1_0 }),
  .out1({ S5718 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6120_ (
  .in1({ S5718, S5717 }),
  .out1({ S5720 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6121_ (
  .in1({ S5720 }),
  .out1({ S5721 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6122_ (
  .in1({ S5363, new_datapath_addsubunit_in1_1 }),
  .out1({ S5722 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6123_ (
  .in1({ S5497, S5410 }),
  .out1({ S5723 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6124_ (
  .in1({ S5722, S5541 }),
  .out1({ S5724 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6125_ (
  .in1({ S5724, S5723 }),
  .out1({ S5725 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6126_ (
  .in1({ S5725, S5721 }),
  .out1({ new_datapath_shiftunit_2355_A })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6127_ (
  .in1({ S5364, S5957 }),
  .out1({ S5726 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6128_ (
  .in1({ S5349, new_datapath_addsubunit_in1_1 }),
  .out1({ S5727 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6129_ (
  .in1({ S5370, new_datapath_addsubunit_in1_0 }),
  .out1({ S5728 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6130_ (
  .in1({ S5442, S5369 }),
  .out1({ S5730 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6131_ (
  .in1({ S5727, S5509 }),
  .out1({ S5731 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6132_ (
  .in1({ S5731, S5726 }),
  .out1({ S5732 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6133_ (
  .in1({ S5728, S5570 }),
  .out1({ S5733 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6134_ (
  .in1({ S5733, S5730 }),
  .out1({ S5734 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6135_ (
  .in1({ S5734, S5732 }),
  .out1({ new_datapath_shiftunit_2373_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6136_ (
  .in1({ S5490, S5411 }),
  .out1({ S5735 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6137_ (
  .in1({ S5591, S5560 }),
  .out1({ S5736 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6138_ (
  .in1({ S5736, S5735 }),
  .out1({ S5737 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6139_ (
  .in1({ S5370, new_datapath_addsubunit_in1_1 }),
  .out1({ S5738 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6140_ (
  .in1({ S5363, new_datapath_addsubunit_in1_3 }),
  .out1({ S5740 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6141_ (
  .in1({ S5740, S5738 }),
  .out1({ S5741 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6142_ (
  .in1({ S5336, new_datapath_addsubunit_in1_0 }),
  .out1({ S5742 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6143_ (
  .in1({ S5349, new_datapath_addsubunit_in1_2 }),
  .out1({ S5743 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6144_ (
  .in1({ S5743, S5742 }),
  .out1({ S5744 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6145_ (
  .in1({ S5744, S5741 }),
  .out1({ S5745 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6146_ (
  .in1({ S5745, S5737 }),
  .out1({ new_datapath_shiftunit_2391_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6147_ (
  .in1({ S5349, new_datapath_addsubunit_in1_3 }),
  .out1({ S5746 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6148_ (
  .in1({ S5370, new_datapath_addsubunit_in1_2 }),
  .out1({ S5747 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6149_ (
  .in1({ S5329, S5975 }),
  .out1({ S5748 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6150_ (
  .in1({ S5336, new_datapath_addsubunit_in1_1 }),
  .out1({ S5750 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6151_ (
  .in1({ S5747, S5746 }),
  .out1({ S5751 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6152_ (
  .in1({ S5580, S5517 }),
  .out1({ S5752 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6153_ (
  .in1({ S5752, S5750 }),
  .out1({ S5753 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6154_ (
  .in1({ S5753, S5751 }),
  .out1({ S5754 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6155_ (
  .in1({ S5616, S5453 }),
  .out1({ S5755 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6156_ (
  .in1({ S5755 }),
  .out1({ S5756 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6157_ (
  .in1({ S5756, S5366 }),
  .out1({ S5757 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6158_ (
  .in1({ S5757, S5748 }),
  .out1({ S5758 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6159_ (
  .in1({ S5758, S5754 }),
  .out1({ new_datapath_shiftunit_2409_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6160_ (
  .in1({ S5370, new_datapath_addsubunit_in1_3 }),
  .out1({ S5760 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6161_ (
  .in1({ S5349, new_datapath_addsubunit_in1_4 }),
  .out1({ S5761 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6162_ (
  .in1({ S5761, S5760 }),
  .out1({ S5762 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6163_ (
  .in1({ S5336, new_datapath_addsubunit_in1_2 }),
  .out1({ S5763 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6164_ (
  .in1({ S5346, new_datapath_addsubunit_in1_0 }),
  .out1({ S5764 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6165_ (
  .in1({ S5764, S5763 }),
  .out1({ S5765 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6166_ (
  .in1({ S5765, S5762 }),
  .out1({ S5766 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6167_ (
  .in1({ S5645, S5601 }),
  .out1({ S5767 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6168_ (
  .in1({ S5477, S5400 }),
  .out1({ S5768 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6169_ (
  .in1({ S5328, new_datapath_addsubunit_in1_1 }),
  .out1({ S5769 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6170_ (
  .in1({ S5769, S5543 }),
  .out1({ S5771 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6171_ (
  .in1({ S5771, S5768 }),
  .out1({ S5772 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6172_ (
  .in1({ S5772 }),
  .out1({ S5773 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6173_ (
  .in1({ S5773, S5767 }),
  .out1({ S5774 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6174_ (
  .in1({ S5774, S5766 }),
  .out1({ new_datapath_shiftunit_2427_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6175_ (
  .in1({ S5336, new_datapath_addsubunit_in1_3 }),
  .out1({ S5775 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6176_ (
  .in1({ S5328, new_datapath_addsubunit_in1_2 }),
  .out1({ S5776 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6177_ (
  .in1({ S5375, new_datapath_addsubunit_in1_0 }),
  .out1({ S5777 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6178_ (
  .in1({ S5346, new_datapath_addsubunit_in1_1 }),
  .out1({ S5778 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6179_ (
  .in1({ S5370, new_datapath_addsubunit_in1_4 }),
  .out1({ S5779 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6180_ (
  .in1({ S5659, S5521 }),
  .out1({ S5781 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6181_ (
  .in1({ S5781, S5454 }),
  .out1({ S5782 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6182_ (
  .in1({ S5617, S5574 }),
  .out1({ S5783 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6183_ (
  .in1({ S5775, S5350 }),
  .out1({ S5784 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6184_ (
  .in1({ S5784, S5783 }),
  .out1({ S5785 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6185_ (
  .in1({ S5785, S5782 }),
  .out1({ S5786 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6186_ (
  .in1({ S5786 }),
  .out1({ S5787 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6187_ (
  .in1({ S5778, S5777 }),
  .out1({ S5788 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6188_ (
  .in1({ S5779, S5776 }),
  .out1({ S5789 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6189_ (
  .in1({ S5789, S5788 }),
  .out1({ S5790 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6190_ (
  .in1({ S5790, S5787 }),
  .out1({ new_datapath_shiftunit_2445_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6191_ (
  .in1({ S5346, new_datapath_addsubunit_in1_2 }),
  .out1({ S5792 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6192_ (
  .in1({ S5328, new_datapath_addsubunit_in1_3 }),
  .out1({ S5793 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6193_ (
  .in1({ S5353, new_datapath_addsubunit_in1_0 }),
  .out1({ S5794 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6194_ (
  .in1({ S5370, new_datapath_addsubunit_in1_5 }),
  .out1({ S5795 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6195_ (
  .in1({ S5375, new_datapath_addsubunit_in1_1 }),
  .out1({ S5796 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6196_ (
  .in1({ S5336, new_datapath_addsubunit_in1_4 }),
  .out1({ S5797 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6197_ (
  .in1({ S5794, S5647 }),
  .out1({ S5798 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6198_ (
  .in1({ S5796, S5405 }),
  .out1({ S5799 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6199_ (
  .in1({ S5799, S5798 }),
  .out1({ S5800 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6200_ (
  .in1({ S5800 }),
  .out1({ S5801 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6201_ (
  .in1({ S5797, S5538 }),
  .out1({ S5802 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6202_ (
  .in1({ S5802, S5801 }),
  .out1({ S5803 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6203_ (
  .in1({ S5792, S5595 }),
  .out1({ S5804 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6204_ (
  .in1({ S5672, S5476 }),
  .out1({ S5805 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6205_ (
  .in1({ S5795, S5793 }),
  .out1({ S5806 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6206_ (
  .in1({ S5806, S5805 }),
  .out1({ S5807 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6207_ (
  .in1({ S5807 }),
  .out1({ S5808 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6208_ (
  .in1({ S5808, S5804 }),
  .out1({ S5809 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6209_ (
  .in1({ S5809, S5803 }),
  .out1({ new_datapath_shiftunit_2463_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6210_ (
  .in1({ S5679, S5662 }),
  .out1({ S5811 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6211_ (
  .in1({ S5353, new_datapath_addsubunit_in1_1 }),
  .out1({ S5812 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6212_ (
  .in1({ S5328, new_datapath_addsubunit_in1_4 }),
  .out1({ S5813 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6213_ (
  .in1({ S5346, new_datapath_addsubunit_in1_3 }),
  .out1({ S5814 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6214_ (
  .in1({ S5337, S5926 }),
  .out1({ S5815 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6215_ (
  .in1({ S5360, new_datapath_addsubunit_in1_0 }),
  .out1({ S5816 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6216_ (
  .in1({ S5375, new_datapath_addsubunit_in1_2 }),
  .out1({ S5817 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6217_ (
  .in1({ S5512, S5445 }),
  .out1({ S5818 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6218_ (
  .in1({ S5818, S5815 }),
  .out1({ S5819 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6219_ (
  .in1({ S5817, S5814 }),
  .out1({ S5820 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6220_ (
  .in1({ S5816, S5813 }),
  .out1({ S5822 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6221_ (
  .in1({ S5822, S5820 }),
  .out1({ S5823 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6222_ (
  .in1({ S5823, S5819 }),
  .out1({ S5824 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6223_ (
  .in1({ S5824 }),
  .out1({ S5825 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6224_ (
  .in1({ S5812, S5625 }),
  .out1({ S5826 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6225_ (
  .in1({ S5826, S5811 }),
  .out1({ S5827 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6226_ (
  .in1({ S5827 }),
  .out1({ S5828 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6227_ (
  .in1({ S5577, S5371 }),
  .out1({ S5829 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6228_ (
  .in1({ S5829, S5828 }),
  .out1({ S5830 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6229_ (
  .in1({ S5830, S5825 }),
  .out1({ new_datapath_shiftunit_2481_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6230_ (
  .in1({ S5353, new_datapath_addsubunit_in1_2 }),
  .out1({ S5831 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6231_ (
  .in1({ S5346, new_datapath_addsubunit_in1_4 }),
  .out1({ S5832 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6232_ (
  .in1({ S5360, new_datapath_addsubunit_in1_1 }),
  .out1({ S5833 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6233_ (
  .in1({ S5328, new_datapath_addsubunit_in1_5 }),
  .out1({ S5834 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6234_ (
  .in1({ S5336, new_datapath_addsubunit_in1_6 }),
  .out1({ S5835 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6235_ (
  .in1({ S5344, new_datapath_addsubunit_in1_0 }),
  .out1({ S5836 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6236_ (
  .in1({ S5375, new_datapath_addsubunit_in1_3 }),
  .out1({ S5837 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6237_ (
  .in1({ S5836, S5833 }),
  .out1({ S5838 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6238_ (
  .in1({ S5834, S5599 }),
  .out1({ S5839 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6239_ (
  .in1({ S5839, S5838 }),
  .out1({ S5840 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6240_ (
  .in1({ S5840 }),
  .out1({ S5842 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6241_ (
  .in1({ S5835, S5675 }),
  .out1({ S5843 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6242_ (
  .in1({ S5843, S5842 }),
  .out1({ S5844 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6243_ (
  .in1({ S5831, S5692 }),
  .out1({ S5845 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6244_ (
  .in1({ S5542, S5489 }),
  .out1({ S5846 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6245_ (
  .in1({ S5846, S5845 }),
  .out1({ S5847 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6246_ (
  .in1({ S5837, S5404 }),
  .out1({ S5848 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6247_ (
  .in1({ S5832, S5634 }),
  .out1({ S5849 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6248_ (
  .in1({ S5849, S5848 }),
  .out1({ S5850 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6249_ (
  .in1({ S5850, S5847 }),
  .out1({ S5851 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6250_ (
  .in1({ S5851 }),
  .out1({ S5853 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6251_ (
  .in1({ S5853, S5844 }),
  .out1({ new_datapath_shiftunit_2499_A })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6252_ (
  .in1({ S5446, S5338 }),
  .out1({ S5854 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6253_ (
  .in1({ S5360, new_datapath_addsubunit_in1_2 }),
  .out1({ S5855 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6254_ (
  .in1({ S5358, new_datapath_addsubunit_in1_0 }),
  .out1({ S5856 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6255_ (
  .in1({ S5375, new_datapath_addsubunit_in1_4 }),
  .out1({ S5857 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6256_ (
  .in1({ S5344, new_datapath_addsubunit_in1_1 }),
  .out1({ S5858 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6257_ (
  .in1({ S5353, new_datapath_addsubunit_in1_3 }),
  .out1({ S5859 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6258_ (
  .in1({ S5328, new_datapath_addsubunit_in1_6 }),
  .out1({ S5860 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6259_ (
  .in1({ S5346, new_datapath_addsubunit_in1_5 }),
  .out1({ S5861 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6260_ (
  .in1({ S5657, S5622 }),
  .out1({ S5863 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6261_ (
  .in1({ S5863, S5854 }),
  .out1({ S5864 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6262_ (
  .in1({ S5861, S5857 }),
  .out1({ S5865 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6263_ (
  .in1({ S5859, S5855 }),
  .out1({ S5866 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6264_ (
  .in1({ S5866, S5865 }),
  .out1({ S5867 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6265_ (
  .in1({ S5867, S5864 }),
  .out1({ S5868 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6266_ (
  .in1({ S5860, S5856 }),
  .out1({ S5869 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6267_ (
  .in1({ S5858, S5698 }),
  .out1({ S5870 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6268_ (
  .in1({ S5870, S5869 }),
  .out1({ S5871 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6269_ (
  .in1({ S5686, S5572 }),
  .out1({ S5872 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6270_ (
  .in1({ S5872, S5514 }),
  .out1({ S5873 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6271_ (
  .in1({ S5873, S5871 }),
  .out1({ S5874 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6272_ (
  .in1({ S5874, S5868 }),
  .out1({ S5875 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6273_ (
  .in1({ S5875 }),
  .out1({ new_datapath_shiftunit_2517_A })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6274_ (
  .in1({ S5361, S5947 }),
  .out1({ S5876 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6275_ (
  .in1({ S5358, new_datapath_addsubunit_in1_1 }),
  .out1({ S5877 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6276_ (
  .in1({ S5396, new_datapath_addsubunit_in1_0 }),
  .out1({ S5878 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6277_ (
  .in1({ S5328, new_datapath_addsubunit_in1_7 }),
  .out1({ S5879 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6278_ (
  .in1({ S5375, new_datapath_addsubunit_in1_5 }),
  .out1({ S5880 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6279_ (
  .in1({ S5880 }),
  .out1({ S5881 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6280_ (
  .in1({ S5346, new_datapath_addsubunit_in1_6 }),
  .out1({ S5883 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6281_ (
  .in1({ S5344, new_datapath_addsubunit_in1_2 }),
  .out1({ S5884 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6282_ (
  .in1({ S5353, new_datapath_addsubunit_in1_4 }),
  .out1({ S5885 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6283_ (
  .in1({ S5884, S5596 }),
  .out1({ S5886 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6284_ (
  .in1({ S5886, S5876 }),
  .out1({ S5887 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6285_ (
  .in1({ S5887, S5878 }),
  .out1({ S5888 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6286_ (
  .in1({ S5635, S5406 }),
  .out1({ S5889 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6287_ (
  .in1({ S5889, S5888 }),
  .out1({ S5890 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6288_ (
  .in1({ S5670, S5539 }),
  .out1({ S5891 })
);
notg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) notg_6289_ (
  .in1({ S5891 }),
  .out1({ S5892 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6290_ (
  .in1({ S5892, S5877 }),
  .out1({ S5894 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6291_ (
  .in1({ S5883, S5879 }),
  .out1({ S5895 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6292_ (
  .in1({ S5895, S5881 }),
  .out1({ S5896 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6293_ (
  .in1({ S5703, S5486 }),
  .out1({ S5897 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6294_ (
  .in1({ S5885, S5694 }),
  .out1({ S5898 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6295_ (
  .in1({ S5898, S5897 }),
  .out1({ S5899 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6296_ (
  .in1({ S5899, S5896 }),
  .out1({ S5900 })
);
nor_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nor_n_6297_ (
  .in1({ S5900, S5894 }),
  .out1({ S5901 })
);
nand_n #(
  .n(32'b00000000000000000000000000000010),
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) nand_n_6298_ (
  .in1({ S5901, S5890 }),
  .out1({ new_datapath_shiftunit_2534_A })
);
bufg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) bufg_6299_ (
  .in1({ new_controller_outflag_7 }),
  .out1({ S3 })
);
bufg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) bufg_6300_ (
  .in1({ new_controller_outflag_0 }),
  .out1({ S66 })
);
bufg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) bufg_6301_ (
  .in1({ new_controller_outflag_1 }),
  .out1({ S67 })
);
bufg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) bufg_6302_ (
  .in1({ new_controller_outflag_2 }),
  .out1({ S68 })
);
bufg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) bufg_6303_ (
  .in1({ new_controller_outflag_3 }),
  .out1({ S69 })
);
bufg #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) bufg_6304_ (
  .in1({ new_controller_outflag_6 }),
  .out1({ S72 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6305_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ new_controller_1423_Y_0 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_pstate_0 }),
  .Si({ S6264 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6306_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ new_controller_1423_Y_1 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_pstate_1 }),
  .Si({ S6265 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6307_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S73 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_adr_outreg_0 }),
  .Si({ S6287 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6308_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S74 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_adr_outreg_1 }),
  .Si({ S6219 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6309_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S75 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_adr_outreg_2 }),
  .Si({ S6273 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6310_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S76 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_adr_outreg_3 }),
  .Si({ S6276 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6311_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S77 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_adr_outreg_4 }),
  .Si({ S6271 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6312_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S78 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_adr_outreg_5 }),
  .Si({ S6280 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6313_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S79 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_adr_outreg_6 }),
  .Si({ S6285 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6314_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S80 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_adr_outreg_7 }),
  .Si({ S6275 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6315_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S81 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_adr_outreg_8 }),
  .Si({ S6286 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6316_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S82 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_adr_outreg_9 }),
  .Si({ S6279 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6317_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S83 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_adr_outreg_10 }),
  .Si({ S6281 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6318_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S84 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_adr_outreg_11 }),
  .Si({ S6282 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6319_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S85 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_adr_outreg_12 }),
  .Si({ S6283 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6320_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S86 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_adr_outreg_13 }),
  .Si({ S6284 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6321_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S87 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_adr_outreg_14 }),
  .Si({ S6278 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6322_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S4 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_adr_outreg_15 }),
  .Si({ S6221 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6323_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S66 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_outflag_0 }),
  .Si({ S6277 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6324_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S67 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_outflag_1 }),
  .Si({ S6274 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6325_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S68 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_outflag_2 }),
  .Si({ S6288 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6326_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S69 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_outflag_3 }),
  .Si({ S6218 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6327_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S70 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_407_B_0 }),
  .Si({ S6217 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6328_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S71 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_407_B_2 }),
  .Si({ S6289 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6329_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S72 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_outflag_6 }),
  .Si({ S6272 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6330_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S3 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_outflag_7 }),
  .Si({ S6306 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6331_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S51 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_instruction_0 }),
  .Si({ S6231 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6332_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S52 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_instruction_1 }),
  .Si({ S6296 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6333_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S53 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_instruction_2 }),
  .Si({ S6228 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6334_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S54 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_instruction_3 }),
  .Si({ S6230 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6335_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S55 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_fib_0 }),
  .Si({ S6227 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6336_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S56 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_fib_1 }),
  .Si({ S6225 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6337_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S57 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_fib_2 }),
  .Si({ S6224 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6338_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S58 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_fib_3 }),
  .Si({ S6295 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6339_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S59 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_fib_4 }),
  .Si({ S6294 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6340_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S60 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_234_B_0 }),
  .Si({ S6291 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6341_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S61 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_opcode_2 }),
  .Si({ S6297 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6342_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S62 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_opcode_3 }),
  .Si({ S6220 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6343_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S63 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_opcode_4 }),
  .Si({ S6229 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6344_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S64 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_opcode_5 }),
  .Si({ S6226 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6345_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S65 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_opcode_6 }),
  .Si({ S6292 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6346_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S2 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_controller_opcode_7 }),
  .Si({ S6268 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6347_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S20 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu1_0 }),
  .Si({ S6234 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6348_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S21 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu1_1 }),
  .Si({ S6233 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6349_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S22 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu1_2 }),
  .Si({ S6254 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6350_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S23 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu1_3 }),
  .Si({ S6253 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6351_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S24 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu1_4 }),
  .Si({ S6232 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6352_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S25 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu1_5 }),
  .Si({ S6259 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6353_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S26 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu1_6 }),
  .Si({ S6258 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6354_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S27 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu1_7 }),
  .Si({ S6257 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6355_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S28 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu1_8 }),
  .Si({ S6252 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6356_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S29 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu1_9 }),
  .Si({ S6251 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6357_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S30 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu1_10 }),
  .Si({ S6250 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6358_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S31 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu1_11 }),
  .Si({ S6249 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6359_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S32 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu1_12 }),
  .Si({ S6248 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6360_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S33 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu1_13 }),
  .Si({ S6247 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6361_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S34 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu1_14 }),
  .Si({ S6256 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6362_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S35 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu1_15 }),
  .Si({ S6246 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6363_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S36 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu2_0 }),
  .Si({ S6245 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6364_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S37 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu2_1 }),
  .Si({ S6244 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6365_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S38 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu2_2 }),
  .Si({ S6243 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6366_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S39 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu2_3 }),
  .Si({ S6242 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6367_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S40 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu2_4 }),
  .Si({ S6241 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6368_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S41 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu2_5 }),
  .Si({ S6240 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6369_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S42 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu2_6 }),
  .Si({ S6239 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6370_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S43 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu2_7 }),
  .Si({ S6238 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6371_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S44 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu2_8 }),
  .Si({ S6237 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6372_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S45 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu2_9 }),
  .Si({ S6293 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6373_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S46 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu2_10 }),
  .Si({ S6236 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6374_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S47 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu2_11 }),
  .Si({ S6290 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6375_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S48 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu2_12 }),
  .Si({ S6235 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6376_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S49 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu2_13 }),
  .Si({ S6298 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6377_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S50 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu2_14 }),
  .Si({ S6255 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6378_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S1 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_multdivunit_outmdu2_15 }),
  .Si({ S6222 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6379_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S5 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_muxmem_in2_0 }),
  .Si({ S6301 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6380_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S6 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_muxmem_in2_1 }),
  .Si({ S6266 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6381_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S7 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_muxmem_in2_2 }),
  .Si({ S6267 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6382_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S8 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_muxmem_in2_3 }),
  .Si({ S6263 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6383_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S9 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_muxmem_in2_4 }),
  .Si({ S6270 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6384_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S10 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_muxmem_in2_5 }),
  .Si({ S6223 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6385_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S11 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_muxmem_in2_6 }),
  .Si({ S6304 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6386_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S12 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_muxmem_in2_7 }),
  .Si({ S6269 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6387_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S13 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_muxmem_in2_8 }),
  .Si({ S6305 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6388_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S14 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_muxmem_in2_9 }),
  .Si({ S6302 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6389_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S15 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_muxmem_in2_10 }),
  .Si({ S6262 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6390_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S16 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_muxmem_in2_11 }),
  .Si({ S6261 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6391_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S17 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_muxmem_in2_12 }),
  .Si({ S6299 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6392_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S18 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_muxmem_in2_13 }),
  .Si({ S6303 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6393_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S19 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_muxmem_in2_14 }),
  .Si({ S6260 }),
  .global_reset({ 1'b0 })
);
dff #(
  .tphl(32'b00000000000000000000000000000000),
  .tplh(32'b00000000000000000000000000000000)
) dff_6394_ (
  .C({ new_controller_clk }),
  .CE({ 1'b1 }),
  .CLR({ new_controller_rst }),
  .D({ S0 }),
  .NbarT({ 1'b0 }),
  .PRE({ 1'b0 }),
  .Q({ new_datapath_muxmem_in2_15 }),
  .Si({ S6300 }),
  .global_reset({ 1'b0 })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6395_ (
  .in1({ new_datapath_addrbus_0 }),
  .out1({ addrBus[0] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6396_ (
  .in1({ new_datapath_addrbus_1 }),
  .out1({ addrBus[1] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6397_ (
  .in1({ new_datapath_addrbus_10 }),
  .out1({ addrBus[10] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6398_ (
  .in1({ new_datapath_addrbus_11 }),
  .out1({ addrBus[11] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6399_ (
  .in1({ new_datapath_addrbus_12 }),
  .out1({ addrBus[12] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6400_ (
  .in1({ new_datapath_addrbus_13 }),
  .out1({ addrBus[13] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6401_ (
  .in1({ new_datapath_addrbus_14 }),
  .out1({ addrBus[14] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6402_ (
  .in1({ new_datapath_addrbus_15 }),
  .out1({ addrBus[15] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6403_ (
  .in1({ new_datapath_addrbus_2 }),
  .out1({ addrBus[2] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6404_ (
  .in1({ new_datapath_addrbus_3 }),
  .out1({ addrBus[3] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6405_ (
  .in1({ new_datapath_addrbus_4 }),
  .out1({ addrBus[4] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6406_ (
  .in1({ new_datapath_addrbus_5 }),
  .out1({ addrBus[5] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6407_ (
  .in1({ new_datapath_addrbus_6 }),
  .out1({ addrBus[6] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6408_ (
  .in1({ new_datapath_addrbus_7 }),
  .out1({ addrBus[7] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6409_ (
  .in1({ new_datapath_addrbus_8 }),
  .out1({ addrBus[8] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6410_ (
  .in1({ new_datapath_addrbus_9 }),
  .out1({ addrBus[9] })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6411_ (
  .in1({ clk }),
  .out1({ new_controller_clk })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6412_ (
  .in1({ dataBusIn[0] }),
  .out1({ new_datapath_databusin_0 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6413_ (
  .in1({ dataBusIn[1] }),
  .out1({ new_datapath_databusin_1 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6414_ (
  .in1({ dataBusIn[10] }),
  .out1({ new_datapath_databusin_10 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6415_ (
  .in1({ dataBusIn[11] }),
  .out1({ new_datapath_databusin_11 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6416_ (
  .in1({ dataBusIn[12] }),
  .out1({ new_datapath_databusin_12 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6417_ (
  .in1({ dataBusIn[13] }),
  .out1({ new_datapath_databusin_13 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6418_ (
  .in1({ dataBusIn[14] }),
  .out1({ new_datapath_databusin_14 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6419_ (
  .in1({ dataBusIn[15] }),
  .out1({ new_datapath_databusin_15 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6420_ (
  .in1({ dataBusIn[2] }),
  .out1({ new_datapath_databusin_2 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6421_ (
  .in1({ dataBusIn[3] }),
  .out1({ new_datapath_databusin_3 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6422_ (
  .in1({ dataBusIn[4] }),
  .out1({ new_datapath_databusin_4 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6423_ (
  .in1({ dataBusIn[5] }),
  .out1({ new_datapath_databusin_5 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6424_ (
  .in1({ dataBusIn[6] }),
  .out1({ new_datapath_databusin_6 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6425_ (
  .in1({ dataBusIn[7] }),
  .out1({ new_datapath_databusin_7 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6426_ (
  .in1({ dataBusIn[8] }),
  .out1({ new_datapath_databusin_8 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6427_ (
  .in1({ dataBusIn[9] }),
  .out1({ new_datapath_databusin_9 })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6428_ (
  .in1({ new_datapath_addsubunit_in1_0 }),
  .out1({ dataBusOut[0] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6429_ (
  .in1({ new_datapath_addsubunit_in1_1 }),
  .out1({ dataBusOut[1] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6430_ (
  .in1({ new_datapath_addsubunit_in1_10 }),
  .out1({ dataBusOut[10] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6431_ (
  .in1({ new_datapath_addsubunit_in1_11 }),
  .out1({ dataBusOut[11] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6432_ (
  .in1({ new_datapath_addsubunit_in1_12 }),
  .out1({ dataBusOut[12] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6433_ (
  .in1({ new_datapath_addsubunit_in1_13 }),
  .out1({ dataBusOut[13] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6434_ (
  .in1({ new_datapath_addsubunit_in1_14 }),
  .out1({ dataBusOut[14] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6435_ (
  .in1({ new_datapath_addsubunit_in1_15 }),
  .out1({ dataBusOut[15] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6436_ (
  .in1({ new_datapath_addsubunit_in1_2 }),
  .out1({ dataBusOut[2] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6437_ (
  .in1({ new_datapath_addsubunit_in1_3 }),
  .out1({ dataBusOut[3] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6438_ (
  .in1({ new_datapath_addsubunit_in1_4 }),
  .out1({ dataBusOut[4] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6439_ (
  .in1({ new_datapath_addsubunit_in1_5 }),
  .out1({ dataBusOut[5] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6440_ (
  .in1({ new_datapath_addsubunit_in1_6 }),
  .out1({ dataBusOut[6] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6441_ (
  .in1({ new_datapath_addsubunit_in1_7 }),
  .out1({ dataBusOut[7] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6442_ (
  .in1({ new_datapath_addsubunit_in1_8 }),
  .out1({ dataBusOut[8] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6443_ (
  .in1({ new_datapath_addsubunit_in1_9 }),
  .out1({ dataBusOut[9] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6444_ (
  .in1({ new_datapath_indatatrf_0 }),
  .out1({ inDataTRF[0] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6445_ (
  .in1({ new_datapath_indatatrf_1 }),
  .out1({ inDataTRF[1] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6446_ (
  .in1({ new_datapath_indatatrf_10 }),
  .out1({ inDataTRF[10] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6447_ (
  .in1({ new_datapath_indatatrf_11 }),
  .out1({ inDataTRF[11] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6448_ (
  .in1({ new_datapath_indatatrf_12 }),
  .out1({ inDataTRF[12] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6449_ (
  .in1({ new_datapath_indatatrf_13 }),
  .out1({ inDataTRF[13] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6450_ (
  .in1({ new_datapath_indatatrf_14 }),
  .out1({ inDataTRF[14] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6451_ (
  .in1({ new_datapath_indatatrf_15 }),
  .out1({ inDataTRF[15] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6452_ (
  .in1({ new_datapath_indatatrf_2 }),
  .out1({ inDataTRF[2] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6453_ (
  .in1({ new_datapath_indatatrf_3 }),
  .out1({ inDataTRF[3] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6454_ (
  .in1({ new_datapath_indatatrf_4 }),
  .out1({ inDataTRF[4] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6455_ (
  .in1({ new_datapath_indatatrf_5 }),
  .out1({ inDataTRF[5] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6456_ (
  .in1({ new_datapath_indatatrf_6 }),
  .out1({ inDataTRF[6] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6457_ (
  .in1({ new_datapath_indatatrf_7 }),
  .out1({ inDataTRF[7] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6458_ (
  .in1({ new_datapath_indatatrf_8 }),
  .out1({ inDataTRF[8] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6459_ (
  .in1({ new_datapath_indatatrf_9 }),
  .out1({ inDataTRF[9] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6460_ (
  .in1({ new_datapath_muxrd_outmux_0 }),
  .out1({ outMuxrd[0] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6461_ (
  .in1({ new_datapath_muxrd_outmux_1 }),
  .out1({ outMuxrd[1] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6462_ (
  .in1({ new_datapath_muxrd_outmux_2 }),
  .out1({ outMuxrd[2] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6463_ (
  .in1({ new_datapath_muxrd_outmux_3 }),
  .out1({ outMuxrd[3] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6464_ (
  .in1({ new_datapath_muxrs1_outmux_0 }),
  .out1({ outMuxrs1[0] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6465_ (
  .in1({ new_datapath_muxrs1_outmux_1 }),
  .out1({ outMuxrs1[1] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6466_ (
  .in1({ new_datapath_muxrs1_outmux_2 }),
  .out1({ outMuxrs1[2] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6467_ (
  .in1({ new_datapath_muxrs1_outmux_3 }),
  .out1({ outMuxrs1[3] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6468_ (
  .in1({ new_datapath_muxrs2_outmux_0 }),
  .out1({ outMuxrs2[0] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6469_ (
  .in1({ new_datapath_muxrs2_outmux_1 }),
  .out1({ outMuxrs2[1] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6470_ (
  .in1({ new_datapath_muxrs2_outmux_2 }),
  .out1({ outMuxrs2[2] })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6471_ (
  .in1({ new_datapath_muxrs2_outmux_3 }),
  .out1({ outMuxrs2[3] })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6472_ (
  .in1({ p1TRF[0] }),
  .out1({ new_datapath_p1trf_0 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6473_ (
  .in1({ p1TRF[1] }),
  .out1({ new_datapath_p1trf_1 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6474_ (
  .in1({ p1TRF[10] }),
  .out1({ new_datapath_addsubunit_in1_10 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6475_ (
  .in1({ p1TRF[11] }),
  .out1({ new_datapath_addsubunit_in1_11 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6476_ (
  .in1({ p1TRF[12] }),
  .out1({ new_datapath_addsubunit_in1_12 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6477_ (
  .in1({ p1TRF[13] }),
  .out1({ new_datapath_addsubunit_in1_13 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6478_ (
  .in1({ p1TRF[14] }),
  .out1({ new_datapath_addsubunit_in1_14 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6479_ (
  .in1({ p1TRF[15] }),
  .out1({ new_datapath_addsubunit_in1_15 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6480_ (
  .in1({ p1TRF[2] }),
  .out1({ new_datapath_p1trf_2 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6481_ (
  .in1({ p1TRF[3] }),
  .out1({ new_datapath_p1trf_3 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6482_ (
  .in1({ p1TRF[4] }),
  .out1({ new_datapath_p1trf_4 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6483_ (
  .in1({ p1TRF[5] }),
  .out1({ new_datapath_p1trf_5 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6484_ (
  .in1({ p1TRF[6] }),
  .out1({ new_datapath_p1trf_6 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6485_ (
  .in1({ p1TRF[7] }),
  .out1({ new_datapath_p1trf_7 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6486_ (
  .in1({ p1TRF[8] }),
  .out1({ new_datapath_addsubunit_in1_8 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6487_ (
  .in1({ p1TRF[9] }),
  .out1({ new_datapath_addsubunit_in1_9 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6488_ (
  .in1({ p2TRF[0] }),
  .out1({ new_datapath_p2trf_0 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6489_ (
  .in1({ p2TRF[1] }),
  .out1({ new_datapath_p2trf_1 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6490_ (
  .in1({ p2TRF[10] }),
  .out1({ new_datapath_multdivunit_1697_B_10 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6491_ (
  .in1({ p2TRF[11] }),
  .out1({ new_datapath_multdivunit_1697_B_11 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6492_ (
  .in1({ p2TRF[12] }),
  .out1({ new_datapath_multdivunit_1697_B_12 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6493_ (
  .in1({ p2TRF[13] }),
  .out1({ new_datapath_multdivunit_1697_B_13 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6494_ (
  .in1({ p2TRF[14] }),
  .out1({ new_datapath_multdivunit_1697_B_14 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6495_ (
  .in1({ p2TRF[15] }),
  .out1({ new_datapath_multdivunit_1697_B_15 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6496_ (
  .in1({ p2TRF[2] }),
  .out1({ new_datapath_p2trf_2 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6497_ (
  .in1({ p2TRF[3] }),
  .out1({ new_datapath_p2trf_3 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6498_ (
  .in1({ p2TRF[4] }),
  .out1({ new_datapath_p2trf_4 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6499_ (
  .in1({ p2TRF[5] }),
  .out1({ new_datapath_p2trf_5 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6500_ (
  .in1({ p2TRF[6] }),
  .out1({ new_datapath_p2trf_6 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6501_ (
  .in1({ p2TRF[7] }),
  .out1({ new_datapath_p2trf_7 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6502_ (
  .in1({ p2TRF[8] }),
  .out1({ new_datapath_multdivunit_1697_B_8 })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6503_ (
  .in1({ p2TRF[9] }),
  .out1({ new_datapath_multdivunit_1697_B_9 })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6504_ (
  .in1({ new_controller_1133_S_0 }),
  .out1({ readInst })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6505_ (
  .in1({ S6215 }),
  .out1({ readMM })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6506_ (
  .in1({ readyMEM }),
  .out1({ new_controller_readymem })
);
pin #(
  .n(32'b00000000000000000000000000000001)
) pin_6507_ (
  .in1({ rst }),
  .out1({ new_controller_rst })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6508_ (
  .in1({ S6216 }),
  .out1({ writeMM })
);
pout #(
  .n(32'b00000000000000000000000000000001)
) pout_6509_ (
  .in1({ new_controller_1133_Y }),
  .out1({ writeTRF })
);

endmodule